
module buffer1_WORD_SIZE8_55 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffern_WORD_SIZE8_LENGTH1_1 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;


  buffer1_WORD_SIZE8_55 gen1_0__buffer ( .in(in), .out(out), .clk(clk), 
        .clear(clear) );
endmodule


module buffer1_WORD_SIZE8_54 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_53 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffern_WORD_SIZE8_LENGTH2_1 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;

  wire   [8:15] intermediates;

  buffer1_WORD_SIZE8_54 gen1_0__buffer ( .in(in), .out(intermediates), .clk(
        clk), .clear(clear) );
  buffer1_WORD_SIZE8_53 gen1_1__buffer ( .in(intermediates), .out(out), .clk(
        clk), .clear(clear) );
endmodule


module buffer1_WORD_SIZE8_52 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_51 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_50 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffern_WORD_SIZE8_LENGTH3_1 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;

  wire   [8:23] intermediates;

  buffer1_WORD_SIZE8_52 gen1_0__buffer ( .in(in), .out(intermediates[8:15]), 
        .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_51 gen1_1__buffer ( .in(intermediates[8:15]), .out(
        intermediates[16:23]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_50 gen1_2__buffer ( .in(intermediates[16:23]), .out(out), 
        .clk(clk), .clear(clear) );
endmodule


module buffer1_WORD_SIZE8_49 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_48 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_47 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_46 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffern_WORD_SIZE8_LENGTH4_1 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;

  wire   [8:31] intermediates;

  buffer1_WORD_SIZE8_49 gen1_0__buffer ( .in(in), .out(intermediates[8:15]), 
        .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_48 gen1_1__buffer ( .in(intermediates[8:15]), .out(
        intermediates[16:23]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_47 gen1_2__buffer ( .in(intermediates[16:23]), .out(
        intermediates[24:31]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_46 gen1_3__buffer ( .in(intermediates[24:31]), .out(out), 
        .clk(clk), .clear(clear) );
endmodule


module buffer1_WORD_SIZE8_45 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_44 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_43 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_42 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_41 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffern_WORD_SIZE8_LENGTH5_1 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;

  wire   [8:39] intermediates;

  buffer1_WORD_SIZE8_45 gen1_0__buffer ( .in(in), .out(intermediates[8:15]), 
        .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_44 gen1_1__buffer ( .in(intermediates[8:15]), .out(
        intermediates[16:23]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_43 gen1_2__buffer ( .in(intermediates[16:23]), .out(
        intermediates[24:31]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_42 gen1_3__buffer ( .in(intermediates[24:31]), .out(
        intermediates[32:39]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_41 gen1_4__buffer ( .in(intermediates[32:39]), .out(out), 
        .clk(clk), .clear(clear) );
endmodule


module buffer1_WORD_SIZE8_40 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_39 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_38 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_37 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_36 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_35 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffern_WORD_SIZE8_LENGTH6_1 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;

  wire   [8:47] intermediates;

  buffer1_WORD_SIZE8_40 gen1_0__buffer ( .in(in), .out(intermediates[8:15]), 
        .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_39 gen1_1__buffer ( .in(intermediates[8:15]), .out(
        intermediates[16:23]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_38 gen1_2__buffer ( .in(intermediates[16:23]), .out(
        intermediates[24:31]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_37 gen1_3__buffer ( .in(intermediates[24:31]), .out(
        intermediates[32:39]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_36 gen1_4__buffer ( .in(intermediates[32:39]), .out(
        intermediates[40:47]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_35 gen1_5__buffer ( .in(intermediates[40:47]), .out(out), 
        .clk(clk), .clear(clear) );
endmodule


module buffer1_WORD_SIZE8_34 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_33 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_32 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_31 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_30 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_29 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_28 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffern_WORD_SIZE8_LENGTH7_1 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;

  wire   [8:55] intermediates;

  buffer1_WORD_SIZE8_34 gen1_0__buffer ( .in(in), .out(intermediates[8:15]), 
        .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_33 gen1_1__buffer ( .in(intermediates[8:15]), .out(
        intermediates[16:23]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_32 gen1_2__buffer ( .in(intermediates[16:23]), .out(
        intermediates[24:31]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_31 gen1_3__buffer ( .in(intermediates[24:31]), .out(
        intermediates[32:39]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_30 gen1_4__buffer ( .in(intermediates[32:39]), .out(
        intermediates[40:47]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_29 gen1_5__buffer ( .in(intermediates[40:47]), .out(
        intermediates[48:55]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_28 gen1_6__buffer ( .in(intermediates[48:55]), .out(out), 
        .clk(clk), .clear(clear) );
endmodule


module buffer1_WORD_SIZE8_27 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffern_WORD_SIZE8_LENGTH1_0 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;


  buffer1_WORD_SIZE8_27 gen1_0__buffer ( .in(in), .out(out), .clk(clk), 
        .clear(clear) );
endmodule


module buffer1_WORD_SIZE8_26 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_25 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffern_WORD_SIZE8_LENGTH2_0 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;

  wire   [8:15] intermediates;

  buffer1_WORD_SIZE8_26 gen1_0__buffer ( .in(in), .out(intermediates), .clk(
        clk), .clear(clear) );
  buffer1_WORD_SIZE8_25 gen1_1__buffer ( .in(intermediates), .out(out), .clk(
        clk), .clear(clear) );
endmodule


module buffer1_WORD_SIZE8_24 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_23 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_22 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffern_WORD_SIZE8_LENGTH3_0 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;

  wire   [8:23] intermediates;

  buffer1_WORD_SIZE8_24 gen1_0__buffer ( .in(in), .out(intermediates[8:15]), 
        .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_23 gen1_1__buffer ( .in(intermediates[8:15]), .out(
        intermediates[16:23]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_22 gen1_2__buffer ( .in(intermediates[16:23]), .out(out), 
        .clk(clk), .clear(clear) );
endmodule


module buffer1_WORD_SIZE8_21 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_20 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_19 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_18 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffern_WORD_SIZE8_LENGTH4_0 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;

  wire   [8:31] intermediates;

  buffer1_WORD_SIZE8_21 gen1_0__buffer ( .in(in), .out(intermediates[8:15]), 
        .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_20 gen1_1__buffer ( .in(intermediates[8:15]), .out(
        intermediates[16:23]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_19 gen1_2__buffer ( .in(intermediates[16:23]), .out(
        intermediates[24:31]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_18 gen1_3__buffer ( .in(intermediates[24:31]), .out(out), 
        .clk(clk), .clear(clear) );
endmodule


module buffer1_WORD_SIZE8_17 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_16 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_15 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_14 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_13 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffern_WORD_SIZE8_LENGTH5_0 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;

  wire   [8:39] intermediates;

  buffer1_WORD_SIZE8_17 gen1_0__buffer ( .in(in), .out(intermediates[8:15]), 
        .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_16 gen1_1__buffer ( .in(intermediates[8:15]), .out(
        intermediates[16:23]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_15 gen1_2__buffer ( .in(intermediates[16:23]), .out(
        intermediates[24:31]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_14 gen1_3__buffer ( .in(intermediates[24:31]), .out(
        intermediates[32:39]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_13 gen1_4__buffer ( .in(intermediates[32:39]), .out(out), 
        .clk(clk), .clear(clear) );
endmodule


module buffer1_WORD_SIZE8_12 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_11 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_10 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_9 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_8 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_7 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffern_WORD_SIZE8_LENGTH6_0 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;

  wire   [8:47] intermediates;

  buffer1_WORD_SIZE8_12 gen1_0__buffer ( .in(in), .out(intermediates[8:15]), 
        .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_11 gen1_1__buffer ( .in(intermediates[8:15]), .out(
        intermediates[16:23]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_10 gen1_2__buffer ( .in(intermediates[16:23]), .out(
        intermediates[24:31]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_9 gen1_3__buffer ( .in(intermediates[24:31]), .out(
        intermediates[32:39]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_8 gen1_4__buffer ( .in(intermediates[32:39]), .out(
        intermediates[40:47]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_7 gen1_5__buffer ( .in(intermediates[40:47]), .out(out), 
        .clk(clk), .clear(clear) );
endmodule


module buffer1_WORD_SIZE8_6 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_5 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_4 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_3 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_2 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_1 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffer1_WORD_SIZE8_0 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;
  wire   n1;

  DFFRNQ_X1 out_reg_0_ ( .D(in[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(in[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(in[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(in[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(in[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(in[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(in[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(in[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module buffern_WORD_SIZE8_LENGTH7_0 ( in, out, clk, clear );
  input [0:7] in;
  output [0:7] out;
  input clk, clear;

  wire   [8:55] intermediates;

  buffer1_WORD_SIZE8_6 gen1_0__buffer ( .in(in), .out(intermediates[8:15]), 
        .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_5 gen1_1__buffer ( .in(intermediates[8:15]), .out(
        intermediates[16:23]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_4 gen1_2__buffer ( .in(intermediates[16:23]), .out(
        intermediates[24:31]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_3 gen1_3__buffer ( .in(intermediates[24:31]), .out(
        intermediates[32:39]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_2 gen1_4__buffer ( .in(intermediates[32:39]), .out(
        intermediates[40:47]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_1 gen1_5__buffer ( .in(intermediates[40:47]), .out(
        intermediates[48:55]), .clk(clk), .clear(clear) );
  buffer1_WORD_SIZE8_0 gen1_6__buffer ( .in(intermediates[48:55]), .out(out), 
        .clk(clk), .clear(clear) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_63_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_63_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_63_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  INV_X1 U7 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U8 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  AND2_X1 U10 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U14 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(B[3]), .ZN(n23) );
  INV_X1 U39 ( .I(A[2]), .ZN(n32) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_63_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .I(A[0]), .ZN(n3) );
  AND2_X1 U2 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U3 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U4 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U5 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U6 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U7 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U8 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U9 ( .I(B[22]), .ZN(n2) );
  INV_X1 U10 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U11 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_63 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_63_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_63_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_62_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_62_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_62_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_62_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_62 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n2), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n2), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_62_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_62_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_61_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_61_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_61_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_61_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_61 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2, n3;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n3), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n2), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n3), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n3), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n3), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n3), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n3), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n3), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n3), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n3), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n3), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n3), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n3), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n3), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n3), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n2), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n2), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n2), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n2), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n2), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n2), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_61_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_61_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
  INV_X1 U5 ( .I(clear), .ZN(n3) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_60_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_60_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_60_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_60_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_60 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2, n3;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n3), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n2), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n3), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n3), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n3), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n3), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n3), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n3), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n3), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n3), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n3), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n3), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n3), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n3), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n3), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n2), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n2), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n2), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n2), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n2), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n2), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_60_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_60_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
  INV_X1 U5 ( .I(clear), .ZN(n3) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_59_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_59_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_59_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_59_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_59 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n2), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n2), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_59_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_59_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_58_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_58_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_58_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_58_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_58 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n2), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n2), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_58_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_58_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_57_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_57_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_57_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_57_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_57 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n2), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n2), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_57_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_57_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_56_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_56_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_56_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_56_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_56 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n2), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n2), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_56_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_56_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_55_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_55_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_55_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n27) );
  INV_X1 U33 ( .I(A[0]), .ZN(n26) );
  INV_X1 U34 ( .I(B[6]), .ZN(n28) );
  INV_X1 U35 ( .I(A[1]), .ZN(n25) );
  INV_X1 U36 ( .I(B[5]), .ZN(n29) );
  INV_X1 U37 ( .I(B[4]), .ZN(n30) );
  INV_X1 U38 ( .I(A[2]), .ZN(n24) );
  INV_X1 U39 ( .I(B[3]), .ZN(n31) );
  INV_X1 U40 ( .I(B[2]), .ZN(n32) );
  INV_X1 U41 ( .I(B[1]), .ZN(n33) );
  INV_X1 U42 ( .I(A[3]), .ZN(n23) );
  INV_X1 U43 ( .I(B[0]), .ZN(n34) );
  INV_X1 U44 ( .I(A[4]), .ZN(n22) );
  INV_X1 U45 ( .I(A[5]), .ZN(n21) );
  INV_X1 U46 ( .I(A[6]), .ZN(n20) );
  INV_X1 U47 ( .I(A[7]), .ZN(n19) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n19), .A2(n27), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n19), .A2(n28), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n19), .A2(n29), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n19), .A2(n30), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n19), .A2(n31), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n19), .A2(n32), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n19), .A2(n33), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n19), .A2(n34), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n27), .A2(n20), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n28), .A2(n20), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n29), .A2(n20), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n30), .A2(n20), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n31), .A2(n20), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n32), .A2(n20), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n33), .A2(n20), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n34), .A2(n20), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n27), .A2(n21), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n28), .A2(n21), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n29), .A2(n21), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n30), .A2(n21), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n31), .A2(n21), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n32), .A2(n21), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n33), .A2(n21), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n34), .A2(n21), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n27), .A2(n22), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n28), .A2(n22), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n29), .A2(n22), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n30), .A2(n22), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n31), .A2(n22), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n32), .A2(n22), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n33), .A2(n22), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n34), .A2(n22), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n27), .A2(n23), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n28), .A2(n23), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n29), .A2(n23), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n30), .A2(n23), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n31), .A2(n23), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n32), .A2(n23), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n33), .A2(n23), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n34), .A2(n23), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n27), .A2(n24), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n28), .A2(n24), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n29), .A2(n24), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n30), .A2(n24), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n31), .A2(n24), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n32), .A2(n24), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n33), .A2(n24), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n34), .A2(n24), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n27), .A2(n25), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n28), .A2(n25), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n29), .A2(n25), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n30), .A2(n25), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n31), .A2(n25), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n32), .A2(n25), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n33), .A2(n25), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n34), .A2(n25), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n27), .A2(n26), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n28), .A2(n26), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n29), .A2(n26), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n30), .A2(n26), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n31), .A2(n26), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n32), .A2(n26), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n33), .A2(n26), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n34), .A2(n26), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_55_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_55 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_55_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_55_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_54_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_54_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_54_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_54_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_54 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_54_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_54_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_53_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_53_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_53_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_53_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_53 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_53_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_53_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_52_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_52_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_52_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_52_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_52 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_52_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_52_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_51_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_51_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_51_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_51_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_51 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_51_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_51_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_50_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_50_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_50_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_50_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_50 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_50_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_50_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_49_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_49_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_49_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_49_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_49 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_49_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_49_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_48_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_48_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_48_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_48_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_48 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_48_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_48_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_47_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_47_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_47_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n27) );
  INV_X1 U33 ( .I(A[0]), .ZN(n26) );
  INV_X1 U34 ( .I(B[6]), .ZN(n28) );
  INV_X1 U35 ( .I(A[1]), .ZN(n25) );
  INV_X1 U36 ( .I(B[5]), .ZN(n29) );
  INV_X1 U37 ( .I(B[4]), .ZN(n30) );
  INV_X1 U38 ( .I(A[2]), .ZN(n24) );
  INV_X1 U39 ( .I(B[3]), .ZN(n31) );
  INV_X1 U40 ( .I(B[2]), .ZN(n32) );
  INV_X1 U41 ( .I(B[1]), .ZN(n33) );
  INV_X1 U42 ( .I(A[3]), .ZN(n23) );
  INV_X1 U43 ( .I(B[0]), .ZN(n34) );
  INV_X1 U44 ( .I(A[4]), .ZN(n22) );
  INV_X1 U45 ( .I(A[5]), .ZN(n21) );
  INV_X1 U46 ( .I(A[6]), .ZN(n20) );
  INV_X1 U47 ( .I(A[7]), .ZN(n19) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n19), .A2(n27), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n19), .A2(n28), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n19), .A2(n29), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n19), .A2(n30), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n19), .A2(n31), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n19), .A2(n32), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n19), .A2(n33), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n19), .A2(n34), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n27), .A2(n20), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n28), .A2(n20), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n29), .A2(n20), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n30), .A2(n20), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n31), .A2(n20), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n32), .A2(n20), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n33), .A2(n20), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n34), .A2(n20), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n27), .A2(n21), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n28), .A2(n21), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n29), .A2(n21), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n30), .A2(n21), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n31), .A2(n21), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n32), .A2(n21), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n33), .A2(n21), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n34), .A2(n21), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n27), .A2(n22), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n28), .A2(n22), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n29), .A2(n22), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n30), .A2(n22), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n31), .A2(n22), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n32), .A2(n22), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n33), .A2(n22), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n34), .A2(n22), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n27), .A2(n23), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n28), .A2(n23), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n29), .A2(n23), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n30), .A2(n23), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n31), .A2(n23), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n32), .A2(n23), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n33), .A2(n23), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n34), .A2(n23), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n27), .A2(n24), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n28), .A2(n24), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n29), .A2(n24), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n30), .A2(n24), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n31), .A2(n24), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n32), .A2(n24), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n33), .A2(n24), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n34), .A2(n24), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n27), .A2(n25), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n28), .A2(n25), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n29), .A2(n25), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n30), .A2(n25), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n31), .A2(n25), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n32), .A2(n25), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n33), .A2(n25), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n34), .A2(n25), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n27), .A2(n26), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n28), .A2(n26), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n29), .A2(n26), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n30), .A2(n26), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n31), .A2(n26), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n32), .A2(n26), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n33), .A2(n26), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n34), .A2(n26), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_47_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_47 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_47_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_47_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_46_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_46_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_46_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_46_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_46 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_46_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_46_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_45_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_45_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_45_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_45_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_45 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_45_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_45_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_44_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_44_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_44_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_44_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_44 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_44_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_44_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_43_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_43_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_43_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_43_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_43 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_43_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_43_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_42_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_42_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_42_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_42_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_42 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_42_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_42_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_41_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_41_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_41_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_41_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_41 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_41_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_41_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_40_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_40_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_40_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_40_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_40 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_40_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_40_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_39_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_39_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_39_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n27) );
  INV_X1 U33 ( .I(A[0]), .ZN(n26) );
  INV_X1 U34 ( .I(B[6]), .ZN(n28) );
  INV_X1 U35 ( .I(A[1]), .ZN(n25) );
  INV_X1 U36 ( .I(B[5]), .ZN(n29) );
  INV_X1 U37 ( .I(B[4]), .ZN(n30) );
  INV_X1 U38 ( .I(A[2]), .ZN(n24) );
  INV_X1 U39 ( .I(B[3]), .ZN(n31) );
  INV_X1 U40 ( .I(B[2]), .ZN(n32) );
  INV_X1 U41 ( .I(B[1]), .ZN(n33) );
  INV_X1 U42 ( .I(A[3]), .ZN(n23) );
  INV_X1 U43 ( .I(B[0]), .ZN(n34) );
  INV_X1 U44 ( .I(A[4]), .ZN(n22) );
  INV_X1 U45 ( .I(A[5]), .ZN(n21) );
  INV_X1 U46 ( .I(A[6]), .ZN(n20) );
  INV_X1 U47 ( .I(A[7]), .ZN(n19) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n19), .A2(n27), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n19), .A2(n28), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n19), .A2(n29), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n19), .A2(n30), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n19), .A2(n31), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n19), .A2(n32), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n19), .A2(n33), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n19), .A2(n34), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n27), .A2(n20), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n28), .A2(n20), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n29), .A2(n20), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n30), .A2(n20), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n31), .A2(n20), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n32), .A2(n20), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n33), .A2(n20), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n34), .A2(n20), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n27), .A2(n21), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n28), .A2(n21), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n29), .A2(n21), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n30), .A2(n21), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n31), .A2(n21), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n32), .A2(n21), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n33), .A2(n21), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n34), .A2(n21), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n27), .A2(n22), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n28), .A2(n22), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n29), .A2(n22), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n30), .A2(n22), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n31), .A2(n22), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n32), .A2(n22), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n33), .A2(n22), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n34), .A2(n22), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n27), .A2(n23), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n28), .A2(n23), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n29), .A2(n23), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n30), .A2(n23), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n31), .A2(n23), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n32), .A2(n23), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n33), .A2(n23), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n34), .A2(n23), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n27), .A2(n24), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n28), .A2(n24), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n29), .A2(n24), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n30), .A2(n24), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n31), .A2(n24), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n32), .A2(n24), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n33), .A2(n24), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n34), .A2(n24), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n27), .A2(n25), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n28), .A2(n25), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n29), .A2(n25), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n30), .A2(n25), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n31), .A2(n25), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n32), .A2(n25), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n33), .A2(n25), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n34), .A2(n25), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n27), .A2(n26), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n28), .A2(n26), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n29), .A2(n26), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n30), .A2(n26), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n31), .A2(n26), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n32), .A2(n26), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n33), .A2(n26), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n34), .A2(n26), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_39_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_39 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_39_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_39_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_38_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_38_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_38_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_38_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_38 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_38_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_38_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_37_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_37_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_37_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_37_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_37 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_37_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_37_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_36_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_36_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_36_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_36_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_36 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_36_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_36_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_35_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_35_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_35_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_35_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_35 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_35_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_35_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_34_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_34_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_34_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_34_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_34 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_34_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_34_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_33_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_33_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_33_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_33_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_33 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_33_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_33_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_32_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_32_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_32_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_32_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_32 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_32_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_32_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_31_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_31_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_31_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n27) );
  INV_X1 U33 ( .I(A[0]), .ZN(n26) );
  INV_X1 U34 ( .I(B[6]), .ZN(n28) );
  INV_X1 U35 ( .I(A[1]), .ZN(n25) );
  INV_X1 U36 ( .I(B[5]), .ZN(n29) );
  INV_X1 U37 ( .I(B[4]), .ZN(n30) );
  INV_X1 U38 ( .I(A[2]), .ZN(n24) );
  INV_X1 U39 ( .I(B[3]), .ZN(n31) );
  INV_X1 U40 ( .I(B[2]), .ZN(n32) );
  INV_X1 U41 ( .I(B[1]), .ZN(n33) );
  INV_X1 U42 ( .I(A[3]), .ZN(n23) );
  INV_X1 U43 ( .I(B[0]), .ZN(n34) );
  INV_X1 U44 ( .I(A[4]), .ZN(n22) );
  INV_X1 U45 ( .I(A[5]), .ZN(n21) );
  INV_X1 U46 ( .I(A[6]), .ZN(n20) );
  INV_X1 U47 ( .I(A[7]), .ZN(n19) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n19), .A2(n27), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n19), .A2(n28), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n19), .A2(n29), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n19), .A2(n30), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n19), .A2(n31), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n19), .A2(n32), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n19), .A2(n33), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n19), .A2(n34), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n27), .A2(n20), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n28), .A2(n20), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n29), .A2(n20), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n30), .A2(n20), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n31), .A2(n20), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n32), .A2(n20), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n33), .A2(n20), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n34), .A2(n20), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n27), .A2(n21), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n28), .A2(n21), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n29), .A2(n21), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n30), .A2(n21), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n31), .A2(n21), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n32), .A2(n21), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n33), .A2(n21), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n34), .A2(n21), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n27), .A2(n22), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n28), .A2(n22), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n29), .A2(n22), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n30), .A2(n22), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n31), .A2(n22), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n32), .A2(n22), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n33), .A2(n22), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n34), .A2(n22), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n27), .A2(n23), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n28), .A2(n23), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n29), .A2(n23), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n30), .A2(n23), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n31), .A2(n23), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n32), .A2(n23), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n33), .A2(n23), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n34), .A2(n23), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n27), .A2(n24), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n28), .A2(n24), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n29), .A2(n24), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n30), .A2(n24), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n31), .A2(n24), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n32), .A2(n24), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n33), .A2(n24), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n34), .A2(n24), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n27), .A2(n25), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n28), .A2(n25), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n29), .A2(n25), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n30), .A2(n25), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n31), .A2(n25), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n32), .A2(n25), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n33), .A2(n25), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n34), .A2(n25), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n27), .A2(n26), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n28), .A2(n26), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n29), .A2(n26), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n30), .A2(n26), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n31), .A2(n26), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n32), .A2(n26), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n33), .A2(n26), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n34), .A2(n26), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_31_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_31 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_31_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_31_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_30_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_30_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_30_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_30_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_30 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_30_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_30_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_29_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_29_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_29_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_29_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_29 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_29_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_29_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_28_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_28_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_28_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_28_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_28 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_28_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_28_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_27_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_27_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_27_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_27_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_27 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_27_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_27_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_26_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_26_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_26_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_26_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_26 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_26_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_26_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_25_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_25_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_25_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_25_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_25 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_25_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_25_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_24_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_24_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_24_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_24_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_24 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_24_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_24_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_23_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_23_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_23_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n27) );
  INV_X1 U33 ( .I(A[0]), .ZN(n26) );
  INV_X1 U34 ( .I(B[6]), .ZN(n28) );
  INV_X1 U35 ( .I(A[1]), .ZN(n25) );
  INV_X1 U36 ( .I(B[5]), .ZN(n29) );
  INV_X1 U37 ( .I(B[4]), .ZN(n30) );
  INV_X1 U38 ( .I(A[2]), .ZN(n24) );
  INV_X1 U39 ( .I(B[3]), .ZN(n31) );
  INV_X1 U40 ( .I(B[2]), .ZN(n32) );
  INV_X1 U41 ( .I(B[1]), .ZN(n33) );
  INV_X1 U42 ( .I(A[3]), .ZN(n23) );
  INV_X1 U43 ( .I(B[0]), .ZN(n34) );
  INV_X1 U44 ( .I(A[4]), .ZN(n22) );
  INV_X1 U45 ( .I(A[5]), .ZN(n21) );
  INV_X1 U46 ( .I(A[6]), .ZN(n20) );
  INV_X1 U47 ( .I(A[7]), .ZN(n19) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n19), .A2(n27), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n19), .A2(n28), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n19), .A2(n29), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n19), .A2(n30), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n19), .A2(n31), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n19), .A2(n32), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n19), .A2(n33), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n19), .A2(n34), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n27), .A2(n20), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n28), .A2(n20), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n29), .A2(n20), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n30), .A2(n20), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n31), .A2(n20), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n32), .A2(n20), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n33), .A2(n20), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n34), .A2(n20), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n27), .A2(n21), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n28), .A2(n21), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n29), .A2(n21), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n30), .A2(n21), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n31), .A2(n21), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n32), .A2(n21), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n33), .A2(n21), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n34), .A2(n21), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n27), .A2(n22), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n28), .A2(n22), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n29), .A2(n22), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n30), .A2(n22), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n31), .A2(n22), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n32), .A2(n22), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n33), .A2(n22), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n34), .A2(n22), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n27), .A2(n23), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n28), .A2(n23), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n29), .A2(n23), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n30), .A2(n23), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n31), .A2(n23), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n32), .A2(n23), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n33), .A2(n23), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n34), .A2(n23), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n27), .A2(n24), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n28), .A2(n24), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n29), .A2(n24), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n30), .A2(n24), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n31), .A2(n24), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n32), .A2(n24), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n33), .A2(n24), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n34), .A2(n24), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n27), .A2(n25), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n28), .A2(n25), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n29), .A2(n25), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n30), .A2(n25), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n31), .A2(n25), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n32), .A2(n25), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n33), .A2(n25), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n34), .A2(n25), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n27), .A2(n26), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n28), .A2(n26), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n29), .A2(n26), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n30), .A2(n26), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n31), .A2(n26), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n32), .A2(n26), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n33), .A2(n26), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n34), .A2(n26), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_23_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_23 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_23_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_23_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_22_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_22_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_22_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_22_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_22 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_22_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_22_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_21_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_21_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_21_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_21_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_21 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_21_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_21_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_20_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_20_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_20_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_20_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_20 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_20_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_20_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_19_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_19_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_19_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_19_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_19 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_19_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_19_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_18_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_18_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_18_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_18_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_18 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1, n2;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n2), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n2), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n2), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n2), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n2), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n2), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n2), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n2), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n2), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n2), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n2), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n2), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n2), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n2), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n2), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n2), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n2), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n2), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n2), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n2), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_18_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_18_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
  INV_X1 U4 ( .I(clear), .ZN(n2) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_17_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_17_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_17_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_17_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_17 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_17_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_17_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_16_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_16_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_16_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_16_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_16 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_16_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_16_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_15_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_15_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_15_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n27) );
  INV_X1 U33 ( .I(A[0]), .ZN(n26) );
  INV_X1 U34 ( .I(B[6]), .ZN(n28) );
  INV_X1 U35 ( .I(A[1]), .ZN(n25) );
  INV_X1 U36 ( .I(B[5]), .ZN(n29) );
  INV_X1 U37 ( .I(B[4]), .ZN(n30) );
  INV_X1 U38 ( .I(A[2]), .ZN(n24) );
  INV_X1 U39 ( .I(B[3]), .ZN(n31) );
  INV_X1 U40 ( .I(B[2]), .ZN(n32) );
  INV_X1 U41 ( .I(B[1]), .ZN(n33) );
  INV_X1 U42 ( .I(A[3]), .ZN(n23) );
  INV_X1 U43 ( .I(B[0]), .ZN(n34) );
  INV_X1 U44 ( .I(A[4]), .ZN(n22) );
  INV_X1 U45 ( .I(A[5]), .ZN(n21) );
  INV_X1 U46 ( .I(A[6]), .ZN(n20) );
  INV_X1 U47 ( .I(A[7]), .ZN(n19) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n19), .A2(n27), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n19), .A2(n28), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n19), .A2(n29), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n19), .A2(n30), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n19), .A2(n31), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n19), .A2(n32), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n19), .A2(n33), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n19), .A2(n34), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n27), .A2(n20), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n28), .A2(n20), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n29), .A2(n20), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n30), .A2(n20), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n31), .A2(n20), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n32), .A2(n20), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n33), .A2(n20), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n34), .A2(n20), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n27), .A2(n21), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n28), .A2(n21), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n29), .A2(n21), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n30), .A2(n21), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n31), .A2(n21), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n32), .A2(n21), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n33), .A2(n21), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n34), .A2(n21), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n27), .A2(n22), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n28), .A2(n22), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n29), .A2(n22), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n30), .A2(n22), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n31), .A2(n22), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n32), .A2(n22), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n33), .A2(n22), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n34), .A2(n22), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n27), .A2(n23), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n28), .A2(n23), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n29), .A2(n23), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n30), .A2(n23), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n31), .A2(n23), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n32), .A2(n23), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n33), .A2(n23), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n34), .A2(n23), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n27), .A2(n24), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n28), .A2(n24), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n29), .A2(n24), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n30), .A2(n24), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n31), .A2(n24), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n32), .A2(n24), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n33), .A2(n24), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n34), .A2(n24), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n27), .A2(n25), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n28), .A2(n25), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n29), .A2(n25), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n30), .A2(n25), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n31), .A2(n25), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n32), .A2(n25), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n33), .A2(n25), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n34), .A2(n25), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n27), .A2(n26), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n28), .A2(n26), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n29), .A2(n26), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n30), .A2(n26), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n31), .A2(n26), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n32), .A2(n26), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n33), .A2(n26), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n34), .A2(n26), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_15_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_15 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_15_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_15_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_14_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_14_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_14_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_14_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_14 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_14_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_14_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_13_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_13_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_13_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_13_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_13 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_13_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_13_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_12_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_12_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_12_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_12_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_12 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_12_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_12_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_11_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_11_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_11_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_11_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_11 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_11_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_11_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_10_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_10_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_10_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_10_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_10 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_10_DW02_mult_0 mult_23 ( .A(a), .B(b), 
        .TC(1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_10_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, 
        mult_out_10_, mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, 
        mult_out_15_, mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, 
        mult_out_20_, mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), 
        .CI(1'b0), .SUM(adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_9_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_9_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_9_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_9_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_9 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_9_DW02_mult_0 mult_23 ( .A(a), .B(b), .TC(
        1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, mult_out_11_, 
        mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, mult_out_16_, 
        mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, mult_out_21_, 
        mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_9_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), .CI(1'b0), .SUM(
        adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_8_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_8_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_8_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_8_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_8 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_8_DW02_mult_0 mult_23 ( .A(a), .B(b), .TC(
        1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, mult_out_11_, 
        mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, mult_out_16_, 
        mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, mult_out_21_, 
        mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_8_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), .CI(1'b0), .SUM(
        adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_7_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_7_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_7_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n27) );
  INV_X1 U33 ( .I(A[0]), .ZN(n26) );
  INV_X1 U34 ( .I(B[6]), .ZN(n28) );
  INV_X1 U35 ( .I(A[1]), .ZN(n25) );
  INV_X1 U36 ( .I(B[5]), .ZN(n29) );
  INV_X1 U37 ( .I(B[4]), .ZN(n30) );
  INV_X1 U38 ( .I(A[2]), .ZN(n24) );
  INV_X1 U39 ( .I(B[3]), .ZN(n31) );
  INV_X1 U40 ( .I(B[2]), .ZN(n32) );
  INV_X1 U41 ( .I(B[1]), .ZN(n33) );
  INV_X1 U42 ( .I(A[3]), .ZN(n23) );
  INV_X1 U43 ( .I(B[0]), .ZN(n34) );
  INV_X1 U44 ( .I(A[4]), .ZN(n22) );
  INV_X1 U45 ( .I(A[5]), .ZN(n21) );
  INV_X1 U46 ( .I(A[6]), .ZN(n20) );
  INV_X1 U47 ( .I(A[7]), .ZN(n19) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n19), .A2(n27), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n19), .A2(n28), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n19), .A2(n29), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n19), .A2(n30), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n19), .A2(n31), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n19), .A2(n32), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n19), .A2(n33), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n19), .A2(n34), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n27), .A2(n20), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n28), .A2(n20), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n29), .A2(n20), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n30), .A2(n20), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n31), .A2(n20), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n32), .A2(n20), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n33), .A2(n20), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n34), .A2(n20), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n27), .A2(n21), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n28), .A2(n21), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n29), .A2(n21), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n30), .A2(n21), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n31), .A2(n21), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n32), .A2(n21), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n33), .A2(n21), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n34), .A2(n21), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n27), .A2(n22), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n28), .A2(n22), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n29), .A2(n22), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n30), .A2(n22), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n31), .A2(n22), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n32), .A2(n22), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n33), .A2(n22), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n34), .A2(n22), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n27), .A2(n23), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n28), .A2(n23), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n29), .A2(n23), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n30), .A2(n23), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n31), .A2(n23), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n32), .A2(n23), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n33), .A2(n23), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n34), .A2(n23), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n27), .A2(n24), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n28), .A2(n24), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n29), .A2(n24), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n30), .A2(n24), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n31), .A2(n24), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n32), .A2(n24), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n33), .A2(n24), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n34), .A2(n24), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n27), .A2(n25), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n28), .A2(n25), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n29), .A2(n25), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n30), .A2(n25), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n31), .A2(n25), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n32), .A2(n25), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n33), .A2(n25), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n34), .A2(n25), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n27), .A2(n26), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n28), .A2(n26), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n29), .A2(n26), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n30), .A2(n26), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n31), .A2(n26), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n32), .A2(n26), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n33), .A2(n26), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n34), .A2(n26), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_7_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_7 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_7_DW02_mult_0 mult_23 ( .A(a), .B(b), .TC(
        1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, mult_out_11_, 
        mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, mult_out_16_, 
        mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, mult_out_21_, 
        mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_7_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), .CI(1'b0), .SUM(
        adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_6_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_6_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_6_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_6_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_6 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_6_DW02_mult_0 mult_23 ( .A(a), .B(b), .TC(
        1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, mult_out_11_, 
        mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, mult_out_16_, 
        mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, mult_out_21_, 
        mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_6_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), .CI(1'b0), .SUM(
        adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_5_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_5_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_5_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_5_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_5 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_5_DW02_mult_0 mult_23 ( .A(a), .B(b), .TC(
        1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, mult_out_11_, 
        mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, mult_out_16_, 
        mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, mult_out_21_, 
        mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_5_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), .CI(1'b0), .SUM(
        adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_4_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_4_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_4_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_4_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_4 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_4_DW02_mult_0 mult_23 ( .A(a), .B(b), .TC(
        1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, mult_out_11_, 
        mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, mult_out_16_, 
        mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, mult_out_21_, 
        mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_4_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), .CI(1'b0), .SUM(
        adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_3_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_3_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_3_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_3_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_3 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_3_DW02_mult_0 mult_23 ( .A(a), .B(b), .TC(
        1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, mult_out_11_, 
        mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, mult_out_16_, 
        mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, mult_out_21_, 
        mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_3_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), .CI(1'b0), .SUM(
        adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_2_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_2_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_2_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_2_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_2 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_2_DW02_mult_0 mult_23 ( .A(a), .B(b), .TC(
        1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, mult_out_11_, 
        mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, mult_out_16_, 
        mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, mult_out_21_, 
        mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_2_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), .CI(1'b0), .SUM(
        adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_1_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_1_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_1_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_1_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_1 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_1_DW02_mult_0 mult_23 ( .A(a), .B(b), .TC(
        1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, mult_out_11_, 
        mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, mult_out_16_, 
        mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, mult_out_21_, 
        mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_1_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), .CI(1'b0), .SUM(
        adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV_X1 U2 ( .I(n9), .ZN(n4) );
  INV_X1 U3 ( .I(n21), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A[7]), .A2(B[7]), .ZN(n11) );
  INV_X1 U5 ( .I(n13), .ZN(n5) );
  INV_X1 U6 ( .I(n23), .ZN(n3) );
  INV_X1 U7 ( .I(n15), .ZN(n1) );
  XOR2_X1 U8 ( .A1(n6), .A2(n7), .Z(SUM[9]) );
  NOR2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n7) );
  XOR2_X1 U10 ( .A1(n10), .A2(n11), .Z(SUM[8]) );
  NAND2_X1 U11 ( .A1(n5), .A2(n12), .ZN(n10) );
  XOR2_X1 U12 ( .A1(B[7]), .A2(A[7]), .Z(SUM[7]) );
  XOR2_X1 U13 ( .A1(n14), .A2(B[13]), .Z(SUM[13]) );
  OAI21_X1 U14 ( .A1(n15), .A2(n16), .B(n17), .ZN(n14) );
  XOR2_X1 U15 ( .A1(n18), .A2(n16), .Z(SUM[12]) );
  AOI21_X1 U16 ( .A1(n2), .A2(n19), .B(n20), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n1), .A2(n17), .ZN(n18) );
  NAND2_X1 U18 ( .A1(B[12]), .A2(A[12]), .ZN(n17) );
  NOR2_X1 U19 ( .A1(B[12]), .A2(A[12]), .ZN(n15) );
  XOR2_X1 U20 ( .A1(n19), .A2(n22), .Z(SUM[11]) );
  NOR2_X1 U21 ( .A1(n20), .A2(n21), .ZN(n22) );
  NOR2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n21) );
  AND2_X1 U23 ( .A1(B[11]), .A2(A[11]), .Z(n20) );
  OAI21_X1 U24 ( .A1(n23), .A2(n24), .B(n25), .ZN(n19) );
  XOR2_X1 U25 ( .A1(n26), .A2(n24), .Z(SUM[10]) );
  AOI21_X1 U26 ( .A1(n6), .A2(n4), .B(n8), .ZN(n24) );
  AND2_X1 U27 ( .A1(B[9]), .A2(A[9]), .Z(n8) );
  NOR2_X1 U28 ( .A1(B[9]), .A2(A[9]), .ZN(n9) );
  OAI21_X1 U29 ( .A1(n11), .A2(n13), .B(n12), .ZN(n6) );
  NAND2_X1 U30 ( .A1(B[8]), .A2(A[8]), .ZN(n12) );
  NOR2_X1 U31 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U32 ( .A1(n3), .A2(n25), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NOR2_X1 U34 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_0_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_, CARRYB_7__2_,
         CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_,
         CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_,
         CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__6_, CARRYB_1__5_, CARRYB_1__4_,
         CARRYB_1__3_, CARRYB_1__2_, CARRYB_1__1_, CARRYB_1__0_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_13_, A2_12_, A2_11_,
         A2_10_, A2_9_, A2_8_, A2_7_, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(CARRYB_1__1_), .CI(SUMB_1__2_), .CO(
        CARRYB_2__1_), .S(SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(CARRYB_1__2_), .CI(SUMB_1__3_), .CO(
        CARRYB_2__2_), .S(SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(CARRYB_1__3_), .CI(SUMB_1__4_), .CO(
        CARRYB_2__3_), .S(SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(CARRYB_1__4_), .CI(SUMB_1__5_), .CO(
        CARRYB_2__4_), .S(SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(CARRYB_1__5_), .CI(SUMB_1__6_), .CO(
        CARRYB_2__5_), .S(SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(CARRYB_1__6_), .CI(ab_1__7_), .CO(
        CARRYB_2__6_), .S(SUMB_2__6_) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_0_DW01_add_1 FS_1 ( .A({1'b0, A1_12_, 
        A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, SUMB_7__0_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .B({A2_13_, A2_12_, A2_11_, A2_10_, A2_9_, 
        A2_8_, A2_7_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[15:2]) );
  INV_X1 U2 ( .I(ab_0__6_), .ZN(n16) );
  INV_X1 U3 ( .I(ab_0__7_), .ZN(n18) );
  INV_X1 U4 ( .I(ab_1__5_), .ZN(n15) );
  INV_X1 U5 ( .I(ab_1__6_), .ZN(n17) );
  AND2_X1 U6 ( .A1(SUMB_7__1_), .A2(CARRYB_7__0_), .Z(A2_7_) );
  AND2_X1 U7 ( .A1(SUMB_7__2_), .A2(CARRYB_7__1_), .Z(A2_8_) );
  INV_X1 U8 ( .I(ab_0__5_), .ZN(n14) );
  INV_X1 U9 ( .I(ab_0__4_), .ZN(n12) );
  INV_X1 U10 ( .I(ab_1__4_), .ZN(n13) );
  INV_X1 U11 ( .I(ab_1__3_), .ZN(n11) );
  INV_X1 U12 ( .I(ab_0__3_), .ZN(n10) );
  INV_X1 U13 ( .I(ab_0__2_), .ZN(n8) );
  INV_X1 U14 ( .I(ab_1__2_), .ZN(n9) );
  INV_X1 U15 ( .I(ab_1__1_), .ZN(n7) );
  AND2_X1 U16 ( .A1(SUMB_7__3_), .A2(CARRYB_7__2_), .Z(A2_9_) );
  INV_X1 U17 ( .I(ab_0__1_), .ZN(n6) );
  INV_X1 U18 ( .I(ab_1__0_), .ZN(n5) );
  AND2_X1 U19 ( .A1(SUMB_7__4_), .A2(CARRYB_7__3_), .Z(A2_10_) );
  AND2_X1 U20 ( .A1(SUMB_7__5_), .A2(CARRYB_7__4_), .Z(A2_11_) );
  AND2_X1 U21 ( .A1(SUMB_7__6_), .A2(CARRYB_7__5_), .Z(A2_12_) );
  INV_X1 U22 ( .I(CARRYB_7__6_), .ZN(n4) );
  INV_X1 U23 ( .I(ab_7__7_), .ZN(n3) );
  NOR2_X1 U24 ( .A1(n15), .A2(n16), .ZN(CARRYB_1__5_) );
  NOR2_X1 U25 ( .A1(n17), .A2(n18), .ZN(CARRYB_1__6_) );
  NOR2_X1 U26 ( .A1(n13), .A2(n14), .ZN(CARRYB_1__4_) );
  NOR2_X1 U27 ( .A1(n11), .A2(n12), .ZN(CARRYB_1__3_) );
  NOR2_X1 U28 ( .A1(n9), .A2(n10), .ZN(CARRYB_1__2_) );
  NOR2_X1 U29 ( .A1(n7), .A2(n8), .ZN(CARRYB_1__1_) );
  NOR2_X1 U30 ( .A1(n5), .A2(n6), .ZN(CARRYB_1__0_) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(A2_13_) );
  INV_X1 U32 ( .I(B[7]), .ZN(n19) );
  INV_X1 U33 ( .I(A[0]), .ZN(n34) );
  INV_X1 U34 ( .I(B[6]), .ZN(n20) );
  INV_X1 U35 ( .I(A[1]), .ZN(n33) );
  INV_X1 U36 ( .I(B[5]), .ZN(n21) );
  INV_X1 U37 ( .I(B[4]), .ZN(n22) );
  INV_X1 U38 ( .I(A[2]), .ZN(n32) );
  INV_X1 U39 ( .I(B[3]), .ZN(n23) );
  INV_X1 U40 ( .I(B[2]), .ZN(n24) );
  INV_X1 U41 ( .I(B[1]), .ZN(n25) );
  INV_X1 U42 ( .I(A[3]), .ZN(n31) );
  INV_X1 U43 ( .I(B[0]), .ZN(n26) );
  INV_X1 U44 ( .I(A[4]), .ZN(n30) );
  INV_X1 U45 ( .I(A[5]), .ZN(n29) );
  INV_X1 U46 ( .I(A[6]), .ZN(n28) );
  INV_X1 U47 ( .I(A[7]), .ZN(n27) );
  XOR2_X1 U48 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .Z(A1_6_) );
  XOR2_X1 U49 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .Z(A1_7_) );
  XOR2_X1 U50 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .Z(A1_8_) );
  XOR2_X1 U51 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .Z(A1_9_) );
  XOR2_X1 U52 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .Z(A1_10_) );
  XOR2_X1 U53 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .Z(A1_11_) );
  XOR2_X1 U54 ( .A1(CARRYB_7__6_), .A2(ab_7__7_), .Z(A1_12_) );
  XOR2_X1 U55 ( .A1(ab_1__0_), .A2(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U56 ( .A1(ab_1__1_), .A2(ab_0__2_), .Z(SUMB_1__1_) );
  XOR2_X1 U57 ( .A1(ab_1__2_), .A2(ab_0__3_), .Z(SUMB_1__2_) );
  XOR2_X1 U58 ( .A1(ab_1__3_), .A2(ab_0__4_), .Z(SUMB_1__3_) );
  XOR2_X1 U59 ( .A1(ab_1__4_), .A2(ab_0__5_), .Z(SUMB_1__4_) );
  XOR2_X1 U60 ( .A1(ab_1__5_), .A2(ab_0__6_), .Z(SUMB_1__5_) );
  XOR2_X1 U61 ( .A1(ab_1__6_), .A2(ab_0__7_), .Z(SUMB_1__6_) );
  NOR2_X1 U63 ( .A1(n27), .A2(n19), .ZN(ab_7__7_) );
  NOR2_X1 U64 ( .A1(n27), .A2(n20), .ZN(ab_7__6_) );
  NOR2_X1 U65 ( .A1(n27), .A2(n21), .ZN(ab_7__5_) );
  NOR2_X1 U66 ( .A1(n27), .A2(n22), .ZN(ab_7__4_) );
  NOR2_X1 U67 ( .A1(n27), .A2(n23), .ZN(ab_7__3_) );
  NOR2_X1 U68 ( .A1(n27), .A2(n24), .ZN(ab_7__2_) );
  NOR2_X1 U69 ( .A1(n27), .A2(n25), .ZN(ab_7__1_) );
  NOR2_X1 U70 ( .A1(n27), .A2(n26), .ZN(ab_7__0_) );
  NOR2_X1 U71 ( .A1(n19), .A2(n28), .ZN(ab_6__7_) );
  NOR2_X1 U72 ( .A1(n20), .A2(n28), .ZN(ab_6__6_) );
  NOR2_X1 U73 ( .A1(n21), .A2(n28), .ZN(ab_6__5_) );
  NOR2_X1 U74 ( .A1(n22), .A2(n28), .ZN(ab_6__4_) );
  NOR2_X1 U75 ( .A1(n23), .A2(n28), .ZN(ab_6__3_) );
  NOR2_X1 U76 ( .A1(n24), .A2(n28), .ZN(ab_6__2_) );
  NOR2_X1 U77 ( .A1(n25), .A2(n28), .ZN(ab_6__1_) );
  NOR2_X1 U78 ( .A1(n26), .A2(n28), .ZN(ab_6__0_) );
  NOR2_X1 U79 ( .A1(n19), .A2(n29), .ZN(ab_5__7_) );
  NOR2_X1 U80 ( .A1(n20), .A2(n29), .ZN(ab_5__6_) );
  NOR2_X1 U81 ( .A1(n21), .A2(n29), .ZN(ab_5__5_) );
  NOR2_X1 U82 ( .A1(n22), .A2(n29), .ZN(ab_5__4_) );
  NOR2_X1 U83 ( .A1(n23), .A2(n29), .ZN(ab_5__3_) );
  NOR2_X1 U84 ( .A1(n24), .A2(n29), .ZN(ab_5__2_) );
  NOR2_X1 U85 ( .A1(n25), .A2(n29), .ZN(ab_5__1_) );
  NOR2_X1 U86 ( .A1(n26), .A2(n29), .ZN(ab_5__0_) );
  NOR2_X1 U87 ( .A1(n19), .A2(n30), .ZN(ab_4__7_) );
  NOR2_X1 U88 ( .A1(n20), .A2(n30), .ZN(ab_4__6_) );
  NOR2_X1 U89 ( .A1(n21), .A2(n30), .ZN(ab_4__5_) );
  NOR2_X1 U90 ( .A1(n22), .A2(n30), .ZN(ab_4__4_) );
  NOR2_X1 U91 ( .A1(n23), .A2(n30), .ZN(ab_4__3_) );
  NOR2_X1 U92 ( .A1(n24), .A2(n30), .ZN(ab_4__2_) );
  NOR2_X1 U93 ( .A1(n25), .A2(n30), .ZN(ab_4__1_) );
  NOR2_X1 U94 ( .A1(n26), .A2(n30), .ZN(ab_4__0_) );
  NOR2_X1 U95 ( .A1(n19), .A2(n31), .ZN(ab_3__7_) );
  NOR2_X1 U96 ( .A1(n20), .A2(n31), .ZN(ab_3__6_) );
  NOR2_X1 U97 ( .A1(n21), .A2(n31), .ZN(ab_3__5_) );
  NOR2_X1 U98 ( .A1(n22), .A2(n31), .ZN(ab_3__4_) );
  NOR2_X1 U99 ( .A1(n23), .A2(n31), .ZN(ab_3__3_) );
  NOR2_X1 U100 ( .A1(n24), .A2(n31), .ZN(ab_3__2_) );
  NOR2_X1 U101 ( .A1(n25), .A2(n31), .ZN(ab_3__1_) );
  NOR2_X1 U102 ( .A1(n26), .A2(n31), .ZN(ab_3__0_) );
  NOR2_X1 U103 ( .A1(n19), .A2(n32), .ZN(ab_2__7_) );
  NOR2_X1 U104 ( .A1(n20), .A2(n32), .ZN(ab_2__6_) );
  NOR2_X1 U105 ( .A1(n21), .A2(n32), .ZN(ab_2__5_) );
  NOR2_X1 U106 ( .A1(n22), .A2(n32), .ZN(ab_2__4_) );
  NOR2_X1 U107 ( .A1(n23), .A2(n32), .ZN(ab_2__3_) );
  NOR2_X1 U108 ( .A1(n24), .A2(n32), .ZN(ab_2__2_) );
  NOR2_X1 U109 ( .A1(n25), .A2(n32), .ZN(ab_2__1_) );
  NOR2_X1 U110 ( .A1(n26), .A2(n32), .ZN(ab_2__0_) );
  NOR2_X1 U111 ( .A1(n19), .A2(n33), .ZN(ab_1__7_) );
  NOR2_X1 U112 ( .A1(n20), .A2(n33), .ZN(ab_1__6_) );
  NOR2_X1 U113 ( .A1(n21), .A2(n33), .ZN(ab_1__5_) );
  NOR2_X1 U114 ( .A1(n22), .A2(n33), .ZN(ab_1__4_) );
  NOR2_X1 U115 ( .A1(n23), .A2(n33), .ZN(ab_1__3_) );
  NOR2_X1 U116 ( .A1(n24), .A2(n33), .ZN(ab_1__2_) );
  NOR2_X1 U117 ( .A1(n25), .A2(n33), .ZN(ab_1__1_) );
  NOR2_X1 U118 ( .A1(n26), .A2(n33), .ZN(ab_1__0_) );
  NOR2_X1 U119 ( .A1(n19), .A2(n34), .ZN(ab_0__7_) );
  NOR2_X1 U120 ( .A1(n20), .A2(n34), .ZN(ab_0__6_) );
  NOR2_X1 U121 ( .A1(n21), .A2(n34), .ZN(ab_0__5_) );
  NOR2_X1 U122 ( .A1(n22), .A2(n34), .ZN(ab_0__4_) );
  NOR2_X1 U123 ( .A1(n23), .A2(n34), .ZN(ab_0__3_) );
  NOR2_X1 U124 ( .A1(n24), .A2(n34), .ZN(ab_0__2_) );
  NOR2_X1 U125 ( .A1(n25), .A2(n34), .ZN(ab_0__1_) );
  NOR2_X1 U126 ( .A1(n26), .A2(n34), .ZN(PRODUCT[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4;
  wire   [23:1] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(carry[16]), .A2(B[16]), .Z(carry[17]) );
  AND2_X1 U2 ( .A1(carry[17]), .A2(B[17]), .Z(carry[18]) );
  AND2_X1 U3 ( .A1(carry[18]), .A2(B[18]), .Z(carry[19]) );
  AND2_X1 U4 ( .A1(carry[19]), .A2(B[19]), .Z(carry[20]) );
  AND2_X1 U5 ( .A1(carry[20]), .A2(B[20]), .Z(carry[21]) );
  AND2_X1 U6 ( .A1(carry[21]), .A2(B[21]), .Z(carry[22]) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(carry[23]) );
  INV_X1 U8 ( .I(B[22]), .ZN(n2) );
  INV_X1 U9 ( .I(carry[22]), .ZN(n1) );
  NOR2_X1 U10 ( .A1(n3), .A2(n4), .ZN(carry[1]) );
  INV_X1 U11 ( .I(A[0]), .ZN(n3) );
  INV_X1 U12 ( .I(B[0]), .ZN(n4) );
  XOR2_X1 U13 ( .A1(B[23]), .A2(carry[23]), .Z(SUM[23]) );
  XOR2_X1 U14 ( .A1(B[22]), .A2(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U15 ( .A1(B[21]), .A2(carry[21]), .Z(SUM[21]) );
  XOR2_X1 U16 ( .A1(B[20]), .A2(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U17 ( .A1(B[19]), .A2(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U18 ( .A1(B[18]), .A2(carry[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A1(B[17]), .A2(carry[17]), .Z(SUM[17]) );
  XOR2_X1 U20 ( .A1(B[16]), .A2(carry[16]), .Z(SUM[16]) );
  XOR2_X1 U21 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
endmodule


module MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_0 ( a, b, a_fwd, b_fwd, out, clk, 
        clear );
  input [0:7] a;
  input [0:7] b;
  output [0:7] a_fwd;
  output [0:7] b_fwd;
  output [0:23] out;
  input clk, clear;
  wire   mult_out_9_, mult_out_8_, mult_out_23_, mult_out_22_, mult_out_21_,
         mult_out_20_, mult_out_19_, mult_out_18_, mult_out_17_, mult_out_16_,
         mult_out_15_, mult_out_14_, mult_out_13_, mult_out_12_, mult_out_11_,
         mult_out_10_, n1;
  wire   [0:23] adder_out;

  DFFRNQ_X1 out_reg_0_ ( .D(adder_out[0]), .CLK(clk), .RN(n1), .Q(out[0]) );
  DFFRNQ_X1 out_reg_1_ ( .D(adder_out[1]), .CLK(clk), .RN(n1), .Q(out[1]) );
  DFFRNQ_X1 out_reg_2_ ( .D(adder_out[2]), .CLK(clk), .RN(n1), .Q(out[2]) );
  DFFRNQ_X1 out_reg_3_ ( .D(adder_out[3]), .CLK(clk), .RN(n1), .Q(out[3]) );
  DFFRNQ_X1 out_reg_4_ ( .D(adder_out[4]), .CLK(clk), .RN(n1), .Q(out[4]) );
  DFFRNQ_X1 out_reg_5_ ( .D(adder_out[5]), .CLK(clk), .RN(n1), .Q(out[5]) );
  DFFRNQ_X1 out_reg_6_ ( .D(adder_out[6]), .CLK(clk), .RN(n1), .Q(out[6]) );
  DFFRNQ_X1 out_reg_7_ ( .D(adder_out[7]), .CLK(clk), .RN(n1), .Q(out[7]) );
  DFFRNQ_X1 out_reg_8_ ( .D(adder_out[8]), .CLK(clk), .RN(n1), .Q(out[8]) );
  DFFRNQ_X1 out_reg_9_ ( .D(adder_out[9]), .CLK(clk), .RN(n1), .Q(out[9]) );
  DFFRNQ_X1 out_reg_10_ ( .D(adder_out[10]), .CLK(clk), .RN(n1), .Q(out[10])
         );
  DFFRNQ_X1 out_reg_11_ ( .D(adder_out[11]), .CLK(clk), .RN(n1), .Q(out[11])
         );
  DFFRNQ_X1 out_reg_12_ ( .D(adder_out[12]), .CLK(clk), .RN(n1), .Q(out[12])
         );
  DFFRNQ_X1 out_reg_13_ ( .D(adder_out[13]), .CLK(clk), .RN(n1), .Q(out[13])
         );
  DFFRNQ_X1 out_reg_14_ ( .D(adder_out[14]), .CLK(clk), .RN(n1), .Q(out[14])
         );
  DFFRNQ_X1 out_reg_15_ ( .D(adder_out[15]), .CLK(clk), .RN(n1), .Q(out[15])
         );
  DFFRNQ_X1 out_reg_16_ ( .D(adder_out[16]), .CLK(clk), .RN(n1), .Q(out[16])
         );
  DFFRNQ_X1 out_reg_17_ ( .D(adder_out[17]), .CLK(clk), .RN(n1), .Q(out[17])
         );
  DFFRNQ_X1 out_reg_18_ ( .D(adder_out[18]), .CLK(clk), .RN(n1), .Q(out[18])
         );
  DFFRNQ_X1 out_reg_19_ ( .D(adder_out[19]), .CLK(clk), .RN(n1), .Q(out[19])
         );
  DFFRNQ_X1 out_reg_20_ ( .D(adder_out[20]), .CLK(clk), .RN(n1), .Q(out[20])
         );
  DFFRNQ_X1 out_reg_21_ ( .D(adder_out[21]), .CLK(clk), .RN(n1), .Q(out[21])
         );
  DFFRNQ_X1 out_reg_22_ ( .D(adder_out[22]), .CLK(clk), .RN(n1), .Q(out[22])
         );
  DFFRNQ_X1 out_reg_23_ ( .D(adder_out[23]), .CLK(clk), .RN(n1), .Q(out[23])
         );
  DFFRNQ_X1 a_fwd_reg_0_ ( .D(a[0]), .CLK(clk), .RN(n1), .Q(a_fwd[0]) );
  DFFRNQ_X1 a_fwd_reg_1_ ( .D(a[1]), .CLK(clk), .RN(n1), .Q(a_fwd[1]) );
  DFFRNQ_X1 a_fwd_reg_2_ ( .D(a[2]), .CLK(clk), .RN(n1), .Q(a_fwd[2]) );
  DFFRNQ_X1 a_fwd_reg_3_ ( .D(a[3]), .CLK(clk), .RN(n1), .Q(a_fwd[3]) );
  DFFRNQ_X1 a_fwd_reg_4_ ( .D(a[4]), .CLK(clk), .RN(n1), .Q(a_fwd[4]) );
  DFFRNQ_X1 a_fwd_reg_5_ ( .D(a[5]), .CLK(clk), .RN(n1), .Q(a_fwd[5]) );
  DFFRNQ_X1 a_fwd_reg_6_ ( .D(a[6]), .CLK(clk), .RN(n1), .Q(a_fwd[6]) );
  DFFRNQ_X1 a_fwd_reg_7_ ( .D(a[7]), .CLK(clk), .RN(n1), .Q(a_fwd[7]) );
  DFFRNQ_X1 b_fwd_reg_0_ ( .D(b[0]), .CLK(clk), .RN(n1), .Q(b_fwd[0]) );
  DFFRNQ_X1 b_fwd_reg_1_ ( .D(b[1]), .CLK(clk), .RN(n1), .Q(b_fwd[1]) );
  DFFRNQ_X1 b_fwd_reg_2_ ( .D(b[2]), .CLK(clk), .RN(n1), .Q(b_fwd[2]) );
  DFFRNQ_X1 b_fwd_reg_3_ ( .D(b[3]), .CLK(clk), .RN(n1), .Q(b_fwd[3]) );
  DFFRNQ_X1 b_fwd_reg_4_ ( .D(b[4]), .CLK(clk), .RN(n1), .Q(b_fwd[4]) );
  DFFRNQ_X1 b_fwd_reg_5_ ( .D(b[5]), .CLK(clk), .RN(n1), .Q(b_fwd[5]) );
  DFFRNQ_X1 b_fwd_reg_6_ ( .D(b[6]), .CLK(clk), .RN(n1), .Q(b_fwd[6]) );
  DFFRNQ_X1 b_fwd_reg_7_ ( .D(b[7]), .CLK(clk), .RN(n1), .Q(b_fwd[7]) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_0_DW02_mult_0 mult_23 ( .A(a), .B(b), .TC(
        1'b0), .PRODUCT({mult_out_8_, mult_out_9_, mult_out_10_, mult_out_11_, 
        mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, mult_out_16_, 
        mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, mult_out_21_, 
        mult_out_22_, mult_out_23_}) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_0_DW01_add_0 add_24 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mult_out_8_, mult_out_9_, mult_out_10_, 
        mult_out_11_, mult_out_12_, mult_out_13_, mult_out_14_, mult_out_15_, 
        mult_out_16_, mult_out_17_, mult_out_18_, mult_out_19_, mult_out_20_, 
        mult_out_21_, mult_out_22_, mult_out_23_}), .B(out), .CI(1'b0), .SUM(
        adder_out) );
  INV_X1 U3 ( .I(clear), .ZN(n1) );
endmodule


module systolic_array_DW01_inc_0 ( A, SUM );
  input [23:0] A;
  output [23:0] SUM;

  wire   [23:2] carry;

  HA_X1 U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  HA_X1 U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  HA_X1 U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  HA_X1 U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  HA_X1 U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  HA_X1 U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  HA_X1 U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  HA_X1 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  HA_X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  HA_X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  HA_X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  HA_X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  HA_X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  HA_X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2_X1 U2 ( .A1(carry[23]), .A2(A[23]), .Z(SUM[23]) );
endmodule


module systolic_array ( clk, rst, top_inputs, left_inputs, compute_done, 
        cycles_count, pe_register_vals );
  input [0:63] top_inputs;
  input [0:63] left_inputs;
  output [23:0] cycles_count;
  output [0:1535] pe_register_vals;
  input clk, rst;
  output compute_done;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N30, N31, N32, N33,
         N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47,
         N48, N49, N50, N51, N52, N53, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118,
         SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120,
         SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122,
         SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124,
         SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126,
         SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128;
  wire   [8:511] left_fwd;
  wire   [8:511] top_fwd;

  DFFSNQ_X1 cycles_count_reg_0_ ( .D(N30), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[0]) );
  DFFSNQ_X1 cycles_count_reg_1_ ( .D(N31), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[1]) );
  DFFSNQ_X1 cycles_count_reg_2_ ( .D(N32), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[2]) );
  DFFSNQ_X1 cycles_count_reg_3_ ( .D(N33), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[3]) );
  DFFSNQ_X1 cycles_count_reg_4_ ( .D(N34), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[4]) );
  DFFSNQ_X1 cycles_count_reg_5_ ( .D(N35), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[5]) );
  DFFSNQ_X1 cycles_count_reg_6_ ( .D(N36), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[6]) );
  DFFSNQ_X1 cycles_count_reg_7_ ( .D(N37), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[7]) );
  DFFSNQ_X1 cycles_count_reg_8_ ( .D(N38), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[8]) );
  DFFSNQ_X1 cycles_count_reg_9_ ( .D(N39), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[9]) );
  DFFSNQ_X1 cycles_count_reg_10_ ( .D(N40), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[10]) );
  DFFSNQ_X1 cycles_count_reg_11_ ( .D(N41), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[11]) );
  DFFSNQ_X1 cycles_count_reg_12_ ( .D(N42), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[12]) );
  DFFSNQ_X1 cycles_count_reg_13_ ( .D(N43), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[13]) );
  DFFSNQ_X1 cycles_count_reg_14_ ( .D(N44), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[14]) );
  DFFSNQ_X1 cycles_count_reg_15_ ( .D(N45), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[15]) );
  DFFSNQ_X1 cycles_count_reg_16_ ( .D(N46), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[16]) );
  DFFSNQ_X1 cycles_count_reg_17_ ( .D(N47), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[17]) );
  DFFSNQ_X1 cycles_count_reg_18_ ( .D(N48), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[18]) );
  DFFSNQ_X1 cycles_count_reg_19_ ( .D(N49), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[19]) );
  DFFSNQ_X1 cycles_count_reg_20_ ( .D(N50), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[20]) );
  DFFSNQ_X1 cycles_count_reg_21_ ( .D(N51), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[21]) );
  DFFSNQ_X1 cycles_count_reg_22_ ( .D(N52), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[22]) );
  DFFSNQ_X1 cycles_count_reg_23_ ( .D(N53), .CLK(clk), .SN(1'b1), .Q(
        cycles_count[23]) );
  DFFSNQ_X1 compute_done_reg ( .D(n30), .CLK(clk), .SN(1'b1), .Q(compute_done)
         );
  AND2_X1 U32 ( .A1(N27), .A2(n35), .Z(N53) );
  AND2_X1 U33 ( .A1(N26), .A2(n36), .Z(N52) );
  AND2_X1 U34 ( .A1(N25), .A2(n36), .Z(N51) );
  AND2_X1 U35 ( .A1(N24), .A2(n36), .Z(N50) );
  AND2_X1 U36 ( .A1(N23), .A2(n36), .Z(N49) );
  AND2_X1 U37 ( .A1(N22), .A2(n36), .Z(N48) );
  AND2_X1 U38 ( .A1(N21), .A2(n37), .Z(N47) );
  AND2_X1 U39 ( .A1(N20), .A2(n37), .Z(N46) );
  AND2_X1 U40 ( .A1(N19), .A2(n37), .Z(N45) );
  AND2_X1 U41 ( .A1(N18), .A2(n37), .Z(N44) );
  AND2_X1 U42 ( .A1(N17), .A2(n37), .Z(N43) );
  AND2_X1 U43 ( .A1(N16), .A2(n38), .Z(N42) );
  AND2_X1 U44 ( .A1(N15), .A2(n38), .Z(N41) );
  AND2_X1 U45 ( .A1(N14), .A2(n38), .Z(N40) );
  AND2_X1 U46 ( .A1(N13), .A2(n38), .Z(N39) );
  AND2_X1 U47 ( .A1(N12), .A2(n38), .Z(N38) );
  AND2_X1 U48 ( .A1(N11), .A2(n39), .Z(N37) );
  AND2_X1 U49 ( .A1(N10), .A2(n39), .Z(N36) );
  AND2_X1 U50 ( .A1(N9), .A2(n39), .Z(N35) );
  AND2_X1 U51 ( .A1(N8), .A2(n39), .Z(N34) );
  AND2_X1 U52 ( .A1(N7), .A2(n39), .Z(N33) );
  AND2_X1 U53 ( .A1(N6), .A2(n40), .Z(N32) );
  AND2_X1 U54 ( .A1(N5), .A2(n40), .Z(N31) );
  AND2_X1 U55 ( .A1(N4), .A2(n40), .Z(N30) );
  buffern_WORD_SIZE8_LENGTH1_1 gen1_1__buffer_inst_c ( .in(top_inputs[48:55]), 
        .out(top_fwd[8:15]), .clk(clk), .clear(n34) );
  buffern_WORD_SIZE8_LENGTH2_1 gen1_2__buffer_inst_c ( .in(top_inputs[40:47]), 
        .out(top_fwd[16:23]), .clk(clk), .clear(n34) );
  buffern_WORD_SIZE8_LENGTH3_1 gen1_3__buffer_inst_c ( .in(top_inputs[32:39]), 
        .out(top_fwd[24:31]), .clk(clk), .clear(n34) );
  buffern_WORD_SIZE8_LENGTH4_1 gen1_4__buffer_inst_c ( .in(top_inputs[24:31]), 
        .out(top_fwd[32:39]), .clk(clk), .clear(n31) );
  buffern_WORD_SIZE8_LENGTH5_1 gen1_5__buffer_inst_c ( .in(top_inputs[16:23]), 
        .out(top_fwd[40:47]), .clk(clk), .clear(n31) );
  buffern_WORD_SIZE8_LENGTH6_1 gen1_6__buffer_inst_c ( .in(top_inputs[8:15]), 
        .out(top_fwd[48:55]), .clk(clk), .clear(n31) );
  buffern_WORD_SIZE8_LENGTH7_1 gen1_7__buffer_inst_c ( .in(top_inputs[0:7]), 
        .out(top_fwd[56:63]), .clk(clk), .clear(n31) );
  buffern_WORD_SIZE8_LENGTH1_0 gen2_1__buffer_inst_r ( .in(left_inputs[48:55]), 
        .out(left_fwd[8:15]), .clk(clk), .clear(n34) );
  buffern_WORD_SIZE8_LENGTH2_0 gen2_2__buffer_inst_r ( .in(left_inputs[40:47]), 
        .out(left_fwd[16:23]), .clk(clk), .clear(n34) );
  buffern_WORD_SIZE8_LENGTH3_0 gen2_3__buffer_inst_r ( .in(left_inputs[32:39]), 
        .out(left_fwd[24:31]), .clk(clk), .clear(n34) );
  buffern_WORD_SIZE8_LENGTH4_0 gen2_4__buffer_inst_r ( .in(left_inputs[24:31]), 
        .out(left_fwd[32:39]), .clk(clk), .clear(n31) );
  buffern_WORD_SIZE8_LENGTH5_0 gen2_5__buffer_inst_r ( .in(left_inputs[16:23]), 
        .out(left_fwd[40:47]), .clk(clk), .clear(n31) );
  buffern_WORD_SIZE8_LENGTH6_0 gen2_6__buffer_inst_r ( .in(left_inputs[8:15]), 
        .out(left_fwd[48:55]), .clk(clk), .clear(n31) );
  buffern_WORD_SIZE8_LENGTH7_0 gen2_7__buffer_inst_r ( .in(left_inputs[0:7]), 
        .out(left_fwd[56:63]), .clk(clk), .clear(n31) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_63 gen3_0__gen4_0__mac_inst ( .a(
        left_inputs[56:63]), .b(top_inputs[56:63]), .a_fwd(left_fwd[64:71]), 
        .b_fwd(top_fwd[64:71]), .out(pe_register_vals[0:23]), .clk(clk), 
        .clear(n31) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_62 gen3_0__gen4_1__mac_inst ( .a(
        left_fwd[64:71]), .b(top_fwd[8:15]), .a_fwd(left_fwd[128:135]), 
        .b_fwd(top_fwd[72:79]), .out(pe_register_vals[24:47]), .clk(clk), 
        .clear(n32) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_61 gen3_0__gen4_2__mac_inst ( .a(
        left_fwd[128:135]), .b(top_fwd[16:23]), .a_fwd(left_fwd[192:199]), 
        .b_fwd(top_fwd[80:87]), .out(pe_register_vals[48:71]), .clk(clk), 
        .clear(n34) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_60 gen3_0__gen4_3__mac_inst ( .a(
        left_fwd[192:199]), .b(top_fwd[24:31]), .a_fwd(left_fwd[256:263]), 
        .b_fwd(top_fwd[88:95]), .out(pe_register_vals[72:95]), .clk(clk), 
        .clear(n34) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_59 gen3_0__gen4_4__mac_inst ( .a(
        left_fwd[256:263]), .b(top_fwd[32:39]), .a_fwd(left_fwd[320:327]), 
        .b_fwd(top_fwd[96:103]), .out(pe_register_vals[96:119]), .clk(clk), 
        .clear(n34) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_58 gen3_0__gen4_5__mac_inst ( .a(
        left_fwd[320:327]), .b(top_fwd[40:47]), .a_fwd(left_fwd[384:391]), 
        .b_fwd(top_fwd[104:111]), .out(pe_register_vals[120:143]), .clk(clk), 
        .clear(n34) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_57 gen3_0__gen4_6__mac_inst ( .a(
        left_fwd[384:391]), .b(top_fwd[48:55]), .a_fwd(left_fwd[448:455]), 
        .b_fwd(top_fwd[112:119]), .out(pe_register_vals[144:167]), .clk(clk), 
        .clear(n34) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_56 gen3_0__gen4_7__mac_inst ( .a(
        left_fwd[448:455]), .b(top_fwd[56:63]), .a_fwd({SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8}), .b_fwd(top_fwd[120:127]), .out(
        pe_register_vals[168:191]), .clk(clk), .clear(n34) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_55 gen3_1__gen4_0__mac_inst ( .a(
        left_fwd[8:15]), .b(top_fwd[64:71]), .a_fwd(left_fwd[72:79]), .b_fwd(
        top_fwd[128:135]), .out(pe_register_vals[192:215]), .clk(clk), .clear(
        n34) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_54 gen3_1__gen4_1__mac_inst ( .a(
        left_fwd[72:79]), .b(top_fwd[72:79]), .a_fwd(left_fwd[136:143]), 
        .b_fwd(top_fwd[136:143]), .out(pe_register_vals[216:239]), .clk(clk), 
        .clear(n34) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_53 gen3_1__gen4_2__mac_inst ( .a(
        left_fwd[136:143]), .b(top_fwd[80:87]), .a_fwd(left_fwd[200:207]), 
        .b_fwd(top_fwd[144:151]), .out(pe_register_vals[240:263]), .clk(clk), 
        .clear(n34) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_52 gen3_1__gen4_3__mac_inst ( .a(
        left_fwd[200:207]), .b(top_fwd[88:95]), .a_fwd(left_fwd[264:271]), 
        .b_fwd(top_fwd[152:159]), .out(pe_register_vals[264:287]), .clk(clk), 
        .clear(n34) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_51 gen3_1__gen4_4__mac_inst ( .a(
        left_fwd[264:271]), .b(top_fwd[96:103]), .a_fwd(left_fwd[328:335]), 
        .b_fwd(top_fwd[160:167]), .out(pe_register_vals[288:311]), .clk(clk), 
        .clear(n34) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_50 gen3_1__gen4_5__mac_inst ( .a(
        left_fwd[328:335]), .b(top_fwd[104:111]), .a_fwd(left_fwd[392:399]), 
        .b_fwd(top_fwd[168:175]), .out(pe_register_vals[312:335]), .clk(clk), 
        .clear(n34) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_49 gen3_1__gen4_6__mac_inst ( .a(
        left_fwd[392:399]), .b(top_fwd[112:119]), .a_fwd(left_fwd[456:463]), 
        .b_fwd(top_fwd[176:183]), .out(pe_register_vals[336:359]), .clk(clk), 
        .clear(n33) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_48 gen3_1__gen4_7__mac_inst ( .a(
        left_fwd[456:463]), .b(top_fwd[120:127]), .a_fwd({
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16}), .b_fwd(
        top_fwd[184:191]), .out(pe_register_vals[360:383]), .clk(clk), .clear(
        n33) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_47 gen3_2__gen4_0__mac_inst ( .a(
        left_fwd[16:23]), .b(top_fwd[128:135]), .a_fwd(left_fwd[80:87]), 
        .b_fwd(top_fwd[192:199]), .out(pe_register_vals[384:407]), .clk(clk), 
        .clear(n33) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_46 gen3_2__gen4_1__mac_inst ( .a(
        left_fwd[80:87]), .b(top_fwd[136:143]), .a_fwd(left_fwd[144:151]), 
        .b_fwd(top_fwd[200:207]), .out(pe_register_vals[408:431]), .clk(clk), 
        .clear(n33) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_45 gen3_2__gen4_2__mac_inst ( .a(
        left_fwd[144:151]), .b(top_fwd[144:151]), .a_fwd(left_fwd[208:215]), 
        .b_fwd(top_fwd[208:215]), .out(pe_register_vals[432:455]), .clk(clk), 
        .clear(n33) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_44 gen3_2__gen4_3__mac_inst ( .a(
        left_fwd[208:215]), .b(top_fwd[152:159]), .a_fwd(left_fwd[272:279]), 
        .b_fwd(top_fwd[216:223]), .out(pe_register_vals[456:479]), .clk(clk), 
        .clear(n33) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_43 gen3_2__gen4_4__mac_inst ( .a(
        left_fwd[272:279]), .b(top_fwd[160:167]), .a_fwd(left_fwd[336:343]), 
        .b_fwd(top_fwd[224:231]), .out(pe_register_vals[480:503]), .clk(clk), 
        .clear(n33) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_42 gen3_2__gen4_5__mac_inst ( .a(
        left_fwd[336:343]), .b(top_fwd[168:175]), .a_fwd(left_fwd[400:407]), 
        .b_fwd(top_fwd[232:239]), .out(pe_register_vals[504:527]), .clk(clk), 
        .clear(n33) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_41 gen3_2__gen4_6__mac_inst ( .a(
        left_fwd[400:407]), .b(top_fwd[176:183]), .a_fwd(left_fwd[464:471]), 
        .b_fwd(top_fwd[240:247]), .out(pe_register_vals[528:551]), .clk(clk), 
        .clear(n33) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_40 gen3_2__gen4_7__mac_inst ( .a(
        left_fwd[464:471]), .b(top_fwd[184:191]), .a_fwd({
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24}), .b_fwd(
        top_fwd[248:255]), .out(pe_register_vals[552:575]), .clk(clk), .clear(
        n33) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_39 gen3_3__gen4_0__mac_inst ( .a(
        left_fwd[24:31]), .b(top_fwd[192:199]), .a_fwd(left_fwd[88:95]), 
        .b_fwd(top_fwd[256:263]), .out(pe_register_vals[576:599]), .clk(clk), 
        .clear(n33) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_38 gen3_3__gen4_1__mac_inst ( .a(
        left_fwd[88:95]), .b(top_fwd[200:207]), .a_fwd(left_fwd[152:159]), 
        .b_fwd(top_fwd[264:271]), .out(pe_register_vals[600:623]), .clk(clk), 
        .clear(n33) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_37 gen3_3__gen4_2__mac_inst ( .a(
        left_fwd[152:159]), .b(top_fwd[208:215]), .a_fwd(left_fwd[216:223]), 
        .b_fwd(top_fwd[272:279]), .out(pe_register_vals[624:647]), .clk(clk), 
        .clear(n33) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_36 gen3_3__gen4_3__mac_inst ( .a(
        left_fwd[216:223]), .b(top_fwd[216:223]), .a_fwd(left_fwd[280:287]), 
        .b_fwd(top_fwd[280:287]), .out(pe_register_vals[648:671]), .clk(clk), 
        .clear(n33) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_35 gen3_3__gen4_4__mac_inst ( .a(
        left_fwd[280:287]), .b(top_fwd[224:231]), .a_fwd(left_fwd[344:351]), 
        .b_fwd(top_fwd[288:295]), .out(pe_register_vals[672:695]), .clk(clk), 
        .clear(n33) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_34 gen3_3__gen4_5__mac_inst ( .a(
        left_fwd[344:351]), .b(top_fwd[232:239]), .a_fwd(left_fwd[408:415]), 
        .b_fwd(top_fwd[296:303]), .out(pe_register_vals[696:719]), .clk(clk), 
        .clear(n33) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_33 gen3_3__gen4_6__mac_inst ( .a(
        left_fwd[408:415]), .b(top_fwd[240:247]), .a_fwd(left_fwd[472:479]), 
        .b_fwd(top_fwd[304:311]), .out(pe_register_vals[720:743]), .clk(clk), 
        .clear(n33) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_32 gen3_3__gen4_7__mac_inst ( .a(
        left_fwd[472:479]), .b(top_fwd[248:255]), .a_fwd({
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32}), .b_fwd(
        top_fwd[312:319]), .out(pe_register_vals[744:767]), .clk(clk), .clear(
        n33) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_31 gen3_4__gen4_0__mac_inst ( .a(
        left_fwd[32:39]), .b(top_fwd[256:263]), .a_fwd(left_fwd[96:103]), 
        .b_fwd(top_fwd[320:327]), .out(pe_register_vals[768:791]), .clk(clk), 
        .clear(n33) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_30 gen3_4__gen4_1__mac_inst ( .a(
        left_fwd[96:103]), .b(top_fwd[264:271]), .a_fwd(left_fwd[160:167]), 
        .b_fwd(top_fwd[328:335]), .out(pe_register_vals[792:815]), .clk(clk), 
        .clear(n33) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_29 gen3_4__gen4_2__mac_inst ( .a(
        left_fwd[160:167]), .b(top_fwd[272:279]), .a_fwd(left_fwd[224:231]), 
        .b_fwd(top_fwd[336:343]), .out(pe_register_vals[816:839]), .clk(clk), 
        .clear(n33) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_28 gen3_4__gen4_3__mac_inst ( .a(
        left_fwd[224:231]), .b(top_fwd[280:287]), .a_fwd(left_fwd[288:295]), 
        .b_fwd(top_fwd[344:351]), .out(pe_register_vals[840:863]), .clk(clk), 
        .clear(n32) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_27 gen3_4__gen4_4__mac_inst ( .a(
        left_fwd[288:295]), .b(top_fwd[288:295]), .a_fwd(left_fwd[352:359]), 
        .b_fwd(top_fwd[352:359]), .out(pe_register_vals[864:887]), .clk(clk), 
        .clear(n32) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_26 gen3_4__gen4_5__mac_inst ( .a(
        left_fwd[352:359]), .b(top_fwd[296:303]), .a_fwd(left_fwd[416:423]), 
        .b_fwd(top_fwd[360:367]), .out(pe_register_vals[888:911]), .clk(clk), 
        .clear(n32) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_25 gen3_4__gen4_6__mac_inst ( .a(
        left_fwd[416:423]), .b(top_fwd[304:311]), .a_fwd(left_fwd[480:487]), 
        .b_fwd(top_fwd[368:375]), .out(pe_register_vals[912:935]), .clk(clk), 
        .clear(n32) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_24 gen3_4__gen4_7__mac_inst ( .a(
        left_fwd[480:487]), .b(top_fwd[312:319]), .a_fwd({
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, 
        SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, 
        SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40}), .b_fwd(
        top_fwd[376:383]), .out(pe_register_vals[936:959]), .clk(clk), .clear(
        n32) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_23 gen3_5__gen4_0__mac_inst ( .a(
        left_fwd[40:47]), .b(top_fwd[320:327]), .a_fwd(left_fwd[104:111]), 
        .b_fwd(top_fwd[384:391]), .out(pe_register_vals[960:983]), .clk(clk), 
        .clear(n32) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_22 gen3_5__gen4_1__mac_inst ( .a(
        left_fwd[104:111]), .b(top_fwd[328:335]), .a_fwd(left_fwd[168:175]), 
        .b_fwd(top_fwd[392:399]), .out(pe_register_vals[984:1007]), .clk(clk), 
        .clear(n32) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_21 gen3_5__gen4_2__mac_inst ( .a(
        left_fwd[168:175]), .b(top_fwd[336:343]), .a_fwd(left_fwd[232:239]), 
        .b_fwd(top_fwd[400:407]), .out(pe_register_vals[1008:1031]), .clk(clk), 
        .clear(n32) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_20 gen3_5__gen4_3__mac_inst ( .a(
        left_fwd[232:239]), .b(top_fwd[344:351]), .a_fwd(left_fwd[296:303]), 
        .b_fwd(top_fwd[408:415]), .out(pe_register_vals[1032:1055]), .clk(clk), 
        .clear(n32) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_19 gen3_5__gen4_4__mac_inst ( .a(
        left_fwd[296:303]), .b(top_fwd[352:359]), .a_fwd(left_fwd[360:367]), 
        .b_fwd(top_fwd[416:423]), .out(pe_register_vals[1056:1079]), .clk(clk), 
        .clear(n32) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_18 gen3_5__gen4_5__mac_inst ( .a(
        left_fwd[360:367]), .b(top_fwd[360:367]), .a_fwd(left_fwd[424:431]), 
        .b_fwd(top_fwd[424:431]), .out(pe_register_vals[1080:1103]), .clk(clk), 
        .clear(n32) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_17 gen3_5__gen4_6__mac_inst ( .a(
        left_fwd[424:431]), .b(top_fwd[368:375]), .a_fwd(left_fwd[488:495]), 
        .b_fwd(top_fwd[432:439]), .out(pe_register_vals[1104:1127]), .clk(clk), 
        .clear(n32) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_16 gen3_5__gen4_7__mac_inst ( .a(
        left_fwd[488:495]), .b(top_fwd[376:383]), .a_fwd({
        SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, 
        SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48}), .b_fwd(
        top_fwd[440:447]), .out(pe_register_vals[1128:1151]), .clk(clk), 
        .clear(n32) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_15 gen3_6__gen4_0__mac_inst ( .a(
        left_fwd[48:55]), .b(top_fwd[384:391]), .a_fwd(left_fwd[112:119]), 
        .b_fwd(top_fwd[448:455]), .out(pe_register_vals[1152:1175]), .clk(clk), 
        .clear(n32) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_14 gen3_6__gen4_1__mac_inst ( .a(
        left_fwd[112:119]), .b(top_fwd[392:399]), .a_fwd(left_fwd[176:183]), 
        .b_fwd(top_fwd[456:463]), .out(pe_register_vals[1176:1199]), .clk(clk), 
        .clear(n32) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_13 gen3_6__gen4_2__mac_inst ( .a(
        left_fwd[176:183]), .b(top_fwd[400:407]), .a_fwd(left_fwd[240:247]), 
        .b_fwd(top_fwd[464:471]), .out(pe_register_vals[1200:1223]), .clk(clk), 
        .clear(n32) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_12 gen3_6__gen4_3__mac_inst ( .a(
        left_fwd[240:247]), .b(top_fwd[408:415]), .a_fwd(left_fwd[304:311]), 
        .b_fwd(top_fwd[472:479]), .out(pe_register_vals[1224:1247]), .clk(clk), 
        .clear(n32) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_11 gen3_6__gen4_4__mac_inst ( .a(
        left_fwd[304:311]), .b(top_fwd[416:423]), .a_fwd(left_fwd[368:375]), 
        .b_fwd(top_fwd[480:487]), .out(pe_register_vals[1248:1271]), .clk(clk), 
        .clear(n32) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_10 gen3_6__gen4_5__mac_inst ( .a(
        left_fwd[368:375]), .b(top_fwd[424:431]), .a_fwd(left_fwd[432:439]), 
        .b_fwd(top_fwd[488:495]), .out(pe_register_vals[1272:1295]), .clk(clk), 
        .clear(n32) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_9 gen3_6__gen4_6__mac_inst ( .a(
        left_fwd[432:439]), .b(top_fwd[432:439]), .a_fwd(left_fwd[496:503]), 
        .b_fwd(top_fwd[496:503]), .out(pe_register_vals[1296:1319]), .clk(clk), 
        .clear(n32) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_8 gen3_6__gen4_7__mac_inst ( .a(
        left_fwd[496:503]), .b(top_fwd[440:447]), .a_fwd({
        SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50, 
        SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, 
        SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54, 
        SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56}), .b_fwd(
        top_fwd[504:511]), .out(pe_register_vals[1320:1343]), .clk(clk), 
        .clear(n31) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_7 gen3_7__gen4_0__mac_inst ( .a(
        left_fwd[56:63]), .b(top_fwd[448:455]), .a_fwd(left_fwd[120:127]), 
        .b_fwd({SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58, 
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62, 
        SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64}), .out(
        pe_register_vals[1344:1367]), .clk(clk), .clear(n31) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_6 gen3_7__gen4_1__mac_inst ( .a(
        left_fwd[120:127]), .b(top_fwd[456:463]), .a_fwd(left_fwd[184:191]), 
        .b_fwd({SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66, 
        SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68, 
        SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70, 
        SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72}), .out(
        pe_register_vals[1368:1391]), .clk(clk), .clear(n31) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_5 gen3_7__gen4_2__mac_inst ( .a(
        left_fwd[184:191]), .b(top_fwd[464:471]), .a_fwd(left_fwd[248:255]), 
        .b_fwd({SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74, 
        SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76, 
        SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78, 
        SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80}), .out(
        pe_register_vals[1392:1415]), .clk(clk), .clear(n31) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_4 gen3_7__gen4_3__mac_inst ( .a(
        left_fwd[248:255]), .b(top_fwd[472:479]), .a_fwd(left_fwd[312:319]), 
        .b_fwd({SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82, 
        SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84, 
        SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86, 
        SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88}), .out(
        pe_register_vals[1416:1439]), .clk(clk), .clear(n31) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_3 gen3_7__gen4_4__mac_inst ( .a(
        left_fwd[312:319]), .b(top_fwd[480:487]), .a_fwd(left_fwd[376:383]), 
        .b_fwd({SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90, 
        SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92, 
        SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94, 
        SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96}), .out(
        pe_register_vals[1440:1463]), .clk(clk), .clear(n31) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_2 gen3_7__gen4_5__mac_inst ( .a(
        left_fwd[376:383]), .b(top_fwd[488:495]), .a_fwd(left_fwd[440:447]), 
        .b_fwd({SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98, 
        SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100, 
        SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102, 
        SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104}), .out(
        pe_register_vals[1464:1487]), .clk(clk), .clear(n31) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_1 gen3_7__gen4_6__mac_inst ( .a(
        left_fwd[440:447]), .b(top_fwd[496:503]), .a_fwd(left_fwd[504:511]), 
        .b_fwd({SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106, 
        SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108, 
        SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110, 
        SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112}), .out(
        pe_register_vals[1488:1511]), .clk(clk), .clear(n31) );
  MAC_IN_WORD_SIZE8_OUT_WORD_SIZE24_0 gen3_7__gen4_7__mac_inst ( .a(
        left_fwd[504:511]), .b(top_fwd[504:511]), .a_fwd({
        SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114, 
        SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116, 
        SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118, 
        SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120}), .b_fwd({
        SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122, 
        SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124, 
        SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126, 
        SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128}), .out(
        pe_register_vals[1512:1535]), .clk(clk), .clear(n31) );
  systolic_array_DW01_inc_0 add_108 ( .A(cycles_count), .SUM({N27, N26, N25, 
        N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, 
        N10, N9, N8, N7, N6, N5, N4}) );
  INV_X1 U56 ( .I(n35), .ZN(n34) );
  INV_X1 U57 ( .I(n35), .ZN(n33) );
  BUF_X2 U58 ( .I(n32), .Z(n31) );
  INV_X1 U59 ( .I(n35), .ZN(n32) );
  INV_X1 U60 ( .I(rst), .ZN(n35) );
  NOR2_X1 U61 ( .A1(n34), .A2(n29), .ZN(n30) );
  NOR2_X1 U62 ( .A1(N28), .A2(compute_done), .ZN(n29) );
  INV_X1 U63 ( .I(rst), .ZN(n36) );
  INV_X1 U64 ( .I(rst), .ZN(n37) );
  INV_X1 U65 ( .I(rst), .ZN(n38) );
  INV_X1 U66 ( .I(rst), .ZN(n39) );
  INV_X1 U67 ( .I(rst), .ZN(n40) );
  INV_X1 U68 ( .I(n41), .ZN(n51) );
  AOI21_X1 U69 ( .A1(cycles_count[2]), .A2(cycles_count[1]), .B(
        cycles_count[3]), .ZN(n41) );
  AOI21_X1 U70 ( .A1(cycles_count[4]), .A2(n51), .B(cycles_count[10]), .ZN(n50) );
  NOR3_X1 U71 ( .A1(cycles_count[11]), .A2(cycles_count[13]), .A3(
        cycles_count[12]), .ZN(n49) );
  OR2_X1 U72 ( .A1(cycles_count[15]), .A2(cycles_count[14]), .Z(n42) );
  NOR4_X1 U73 ( .A1(n42), .A2(cycles_count[16]), .A3(cycles_count[18]), .A4(
        cycles_count[17]), .ZN(n48) );
  NOR2_X1 U74 ( .A1(cycles_count[20]), .A2(cycles_count[19]), .ZN(n46) );
  NOR3_X1 U75 ( .A1(cycles_count[21]), .A2(cycles_count[23]), .A3(
        cycles_count[22]), .ZN(n45) );
  NOR2_X1 U76 ( .A1(cycles_count[6]), .A2(cycles_count[5]), .ZN(n44) );
  NOR3_X1 U77 ( .A1(cycles_count[7]), .A2(cycles_count[9]), .A3(
        cycles_count[8]), .ZN(n43) );
  AND4_X1 U78 ( .A1(n46), .A2(n45), .A3(n44), .A4(n43), .Z(n47) );
  NAND4_X1 U79 ( .A1(n50), .A2(n49), .A3(n48), .A4(n47), .ZN(N28) );
endmodule

