# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2014, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *       NGLibraryCreator, Development_version_64 - build 201405300513        *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on us19.nangate.us for user Lucio Rech (lre).
# Local time is now Tue, 3 Jun 2014, 13:07:07.
# Main process id is 12480.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO AND2_X1
  CLASS core ;
  FOREIGN AND2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.256 0.206 0.6959 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.127 0.078 0.525 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.114 0.334 0.64 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.27 0.796 ;
        RECT 0.27 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.162 0.1419 0.19 ;
        RECT 0.114 0.19 0.1419 0.428 ;
        RECT 0.114 0.428 0.1419 0.544 ;
        RECT 0.1419 0.162 0.242 0.19 ;
        RECT 0.242 0.162 0.27 0.19 ;
        RECT 0.242 0.19 0.27 0.428 ;
      LAYER M1 ;
        RECT 0.114 0.162 0.1419 0.19 ;
        RECT 0.114 0.19 0.1419 0.428 ;
        RECT 0.114 0.428 0.1419 0.544 ;
        RECT 0.1419 0.162 0.242 0.19 ;
        RECT 0.242 0.162 0.27 0.19 ;
        RECT 0.242 0.19 0.27 0.428 ;
  END
END AND2_X1

MACRO AND2_X2
  CLASS core ;
  FOREIGN AND2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.448 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.256 0.206 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.248 0.083 0.52 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.302 0.064 0.306 0.13 ;
        RECT 0.302 0.638 0.306 0.704 ;
        RECT 0.306 0.064 0.334 0.13 ;
        RECT 0.306 0.13 0.334 0.638 ;
        RECT 0.306 0.638 0.334 0.704 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.27 0.796 ;
        RECT 0.27 0.74 0.458 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.458 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.054 0.574 0.082 0.602 ;
        RECT 0.082 0.166 0.242 0.194 ;
        RECT 0.082 0.574 0.242 0.602 ;
        RECT 0.242 0.166 0.27 0.194 ;
        RECT 0.242 0.194 0.27 0.574 ;
        RECT 0.242 0.574 0.27 0.602 ;
      LAYER M1 ;
        RECT 0.054 0.574 0.082 0.602 ;
        RECT 0.082 0.166 0.242 0.194 ;
        RECT 0.082 0.574 0.242 0.602 ;
        RECT 0.242 0.166 0.27 0.194 ;
        RECT 0.242 0.194 0.27 0.574 ;
        RECT 0.242 0.574 0.27 0.602 ;
  END
END AND2_X2

MACRO AND3_X1
  CLASS core ;
  FOREIGN AND3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.192 0.334 0.576 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1729 0.192 0.211 0.576 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.048 0.192 0.08 0.576 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.114 0.462 0.654 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.398 0.796 ;
        RECT 0.398 0.74 0.522 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.522 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.079 0.1 0.238 0.132 ;
        RECT 0.054 0.631 0.274 0.659 ;
        RECT 0.274 0.095 0.37 0.137 ;
        RECT 0.274 0.631 0.37 0.659 ;
        RECT 0.37 0.095 0.398 0.137 ;
        RECT 0.37 0.137 0.398 0.631 ;
        RECT 0.37 0.631 0.398 0.659 ;
      LAYER M1 ;
        RECT 0.079 0.1 0.238 0.132 ;
        RECT 0.054 0.631 0.274 0.659 ;
        RECT 0.274 0.095 0.37 0.137 ;
        RECT 0.274 0.631 0.37 0.659 ;
        RECT 0.37 0.095 0.398 0.137 ;
        RECT 0.37 0.137 0.398 0.631 ;
        RECT 0.37 0.631 0.398 0.659 ;
  END
END AND3_X1

MACRO AND3_X2
  CLASS core ;
  FOREIGN AND3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.32 0.206 0.513 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.256 0.083 0.512 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.302 0.27 0.537 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.366 0.064 0.37 0.157 ;
        RECT 0.366 0.638 0.37 0.704 ;
        RECT 0.37 0.064 0.398 0.157 ;
        RECT 0.37 0.157 0.398 0.638 ;
        RECT 0.37 0.638 0.398 0.704 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.334 0.796 ;
        RECT 0.334 0.74 0.522 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.522 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.072 0.08 0.156 ;
        RECT 0.048 0.156 0.08 0.188 ;
        RECT 0.08 0.156 0.298 0.188 ;
        RECT 0.054 0.581 0.146 0.613 ;
        RECT 0.146 0.224 0.306 0.252 ;
        RECT 0.146 0.581 0.306 0.613 ;
        RECT 0.306 0.224 0.334 0.252 ;
        RECT 0.306 0.252 0.334 0.581 ;
        RECT 0.306 0.581 0.334 0.613 ;
      LAYER M1 ;
        RECT 0.048 0.072 0.08 0.156 ;
        RECT 0.048 0.156 0.08 0.188 ;
        RECT 0.08 0.156 0.298 0.188 ;
        RECT 0.054 0.581 0.146 0.613 ;
        RECT 0.146 0.224 0.306 0.252 ;
        RECT 0.146 0.581 0.306 0.613 ;
        RECT 0.306 0.224 0.334 0.252 ;
        RECT 0.306 0.252 0.334 0.581 ;
        RECT 0.306 0.581 0.334 0.613 ;
  END
END AND3_X2

MACRO AND4_X1
  CLASS core ;
  FOREIGN AND4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.192 0.398 0.576 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.24 0.192 0.272 0.576 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.192 0.1419 0.512 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.576 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.114 0.526 0.654 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.462 0.796 ;
        RECT 0.462 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.082 0.636 0.338 0.668 ;
        RECT 0.338 0.1 0.434 0.132 ;
        RECT 0.338 0.636 0.434 0.668 ;
        RECT 0.434 0.1 0.462 0.132 ;
        RECT 0.434 0.132 0.462 0.636 ;
        RECT 0.434 0.636 0.462 0.668 ;
        RECT 0.1409 0.099 0.298 0.147 ;
      LAYER M1 ;
        RECT 0.082 0.636 0.338 0.668 ;
        RECT 0.338 0.1 0.434 0.132 ;
        RECT 0.338 0.636 0.434 0.668 ;
        RECT 0.434 0.1 0.462 0.132 ;
        RECT 0.434 0.132 0.462 0.636 ;
        RECT 0.434 0.636 0.462 0.668 ;
        RECT 0.1409 0.099 0.298 0.147 ;
  END
END AND4_X1

MACRO AND4_X2
  CLASS core ;
  FOREIGN AND4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.64 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.241 0.398 0.576 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.192 0.27 0.577 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.192 0.1419 0.577 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.577 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.096 0.526 0.64 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.462 0.796 ;
        RECT 0.462 0.74 0.65 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.65 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.1419 0.1 0.298 0.132 ;
        RECT 0.082 0.636 0.342 0.668 ;
        RECT 0.342 0.165 0.434 0.197 ;
        RECT 0.342 0.636 0.434 0.668 ;
        RECT 0.434 0.165 0.462 0.197 ;
        RECT 0.434 0.197 0.462 0.636 ;
        RECT 0.434 0.636 0.462 0.668 ;
      LAYER M1 ;
        RECT 0.1419 0.1 0.298 0.132 ;
        RECT 0.082 0.636 0.342 0.668 ;
        RECT 0.342 0.165 0.434 0.197 ;
        RECT 0.342 0.636 0.434 0.668 ;
        RECT 0.434 0.165 0.462 0.197 ;
        RECT 0.434 0.197 0.462 0.636 ;
        RECT 0.434 0.636 0.462 0.668 ;
  END
END AND4_X2

MACRO ANTENNA
  CLASS core ;
  FOREIGN ANTENNA 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.192 BY 0.768 ;
END ANTENNA

MACRO AOI21_X1
  CLASS core ;
  FOREIGN AOI21_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.192 0.206 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.134 0.078 0.512 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.192 0.334 0.512 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.1 0.1419 0.132 ;
        RECT 0.114 0.132 0.1419 0.536 ;
        RECT 0.1419 0.1 0.306 0.132 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.298 0.796 ;
        RECT 0.298 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.58 0.08 0.612 ;
        RECT 0.048 0.612 0.08 0.704 ;
        RECT 0.08 0.58 0.298 0.612 ;
      LAYER M1 ;
        RECT 0.048 0.58 0.08 0.612 ;
        RECT 0.048 0.612 0.08 0.704 ;
        RECT 0.08 0.58 0.298 0.612 ;
  END
END AOI21_X1

MACRO AOI21_X2
  CLASS core ;
  FOREIGN AOI21_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.302 0.398 0.448 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.23 0.27 0.258 ;
        RECT 0.242 0.258 0.27 0.448 ;
        RECT 0.242 0.448 0.27 0.512 ;
        RECT 0.27 0.23 0.493 0.258 ;
        RECT 0.493 0.23 0.531 0.258 ;
        RECT 0.493 0.258 0.531 0.448 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.1419 0.448 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.077 0.166 0.178 0.194 ;
        RECT 0.178 0.166 0.206 0.194 ;
        RECT 0.178 0.194 0.206 0.489 ;
        RECT 0.178 0.489 0.206 0.5709 ;
        RECT 0.178 0.5709 0.206 0.599 ;
        RECT 0.206 0.166 0.43 0.194 ;
        RECT 0.206 0.5709 0.43 0.599 ;
        RECT 0.43 0.5709 0.434 0.599 ;
        RECT 0.434 0.489 0.462 0.5709 ;
        RECT 0.434 0.5709 0.462 0.599 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.526 0.796 ;
        RECT 0.526 0.74 0.535 0.796 ;
        RECT 0.535 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.55 0.08 0.635 ;
        RECT 0.048 0.635 0.08 0.669 ;
        RECT 0.08 0.635 0.498 0.669 ;
        RECT 0.498 0.516 0.526 0.55 ;
        RECT 0.498 0.55 0.526 0.635 ;
        RECT 0.498 0.635 0.526 0.669 ;
        RECT 0.146 0.1019 0.535 0.13 ;
      LAYER M1 ;
        RECT 0.048 0.55 0.08 0.635 ;
        RECT 0.048 0.635 0.08 0.669 ;
        RECT 0.08 0.635 0.498 0.669 ;
        RECT 0.498 0.516 0.526 0.55 ;
        RECT 0.498 0.55 0.526 0.635 ;
        RECT 0.498 0.635 0.526 0.669 ;
        RECT 0.146 0.1019 0.535 0.13 ;
  END
END AOI21_X2

MACRO AOI22_X1
  CLASS core ;
  FOREIGN AOI22_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.448 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.192 0.27 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.192 0.398 0.485 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.198 0.1419 0.576 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.576 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1409 0.1019 0.306 0.13 ;
        RECT 0.306 0.1019 0.334 0.13 ;
        RECT 0.306 0.13 0.334 0.582 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.398 0.796 ;
        RECT 0.398 0.74 0.458 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.458 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.082 0.63 0.37 0.674 ;
        RECT 0.37 0.553 0.398 0.63 ;
        RECT 0.37 0.63 0.398 0.674 ;
      LAYER M1 ;
        RECT 0.082 0.63 0.37 0.674 ;
        RECT 0.37 0.553 0.398 0.63 ;
        RECT 0.37 0.63 0.398 0.674 ;
  END
END AOI22_X1

MACRO AOI22_X2
  CLASS core ;
  FOREIGN AOI22_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.768 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.274 0.462 0.302 ;
        RECT 0.434 0.302 0.462 0.489 ;
        RECT 0.434 0.489 0.462 0.512 ;
        RECT 0.462 0.274 0.654 0.302 ;
        RECT 0.654 0.274 0.6899 0.302 ;
        RECT 0.6899 0.274 0.718 0.302 ;
        RECT 0.6899 0.302 0.718 0.489 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.562 0.37 0.59 0.512 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.306 0.334 0.526 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.242 0.078 0.512 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.2 0.27 0.228 ;
        RECT 0.242 0.228 0.27 0.229 ;
        RECT 0.242 0.229 0.27 0.32 ;
        RECT 0.27 0.2 0.362 0.228 ;
        RECT 0.362 0.2 0.37 0.228 ;
        RECT 0.37 0.2 0.398 0.228 ;
        RECT 0.37 0.228 0.398 0.229 ;
        RECT 0.37 0.229 0.398 0.32 ;
        RECT 0.37 0.32 0.398 0.463 ;
        RECT 0.37 0.463 0.398 0.5679 ;
        RECT 0.37 0.5679 0.398 0.602 ;
        RECT 0.398 0.2 0.626 0.228 ;
        RECT 0.398 0.228 0.626 0.229 ;
        RECT 0.398 0.5679 0.626 0.602 ;
        RECT 0.626 0.2 0.654 0.228 ;
        RECT 0.626 0.228 0.654 0.229 ;
        RECT 0.626 0.463 0.654 0.5679 ;
        RECT 0.626 0.5679 0.654 0.602 ;
        RECT 0.654 0.2 0.6899 0.228 ;
        RECT 0.654 0.228 0.6899 0.229 ;
        RECT 0.6899 0.096 0.718 0.2 ;
        RECT 0.6899 0.2 0.718 0.228 ;
        RECT 0.6899 0.228 0.718 0.229 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.718 0.796 ;
        RECT 0.718 0.74 0.778 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.778 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.406 0.132 0.626 0.164 ;
        RECT 0.626 0.072 0.654 0.132 ;
        RECT 0.626 0.132 0.654 0.164 ;
        RECT 0.077 0.638 0.6899 0.666 ;
        RECT 0.6899 0.557 0.718 0.638 ;
        RECT 0.6899 0.638 0.718 0.666 ;
        RECT 0.0859 0.0869 0.362 0.145 ;
      LAYER M1 ;
        RECT 0.406 0.132 0.626 0.164 ;
        RECT 0.626 0.072 0.654 0.132 ;
        RECT 0.626 0.132 0.654 0.164 ;
        RECT 0.077 0.638 0.6899 0.666 ;
        RECT 0.6899 0.557 0.718 0.638 ;
        RECT 0.6899 0.638 0.718 0.666 ;
        RECT 0.0859 0.0869 0.362 0.145 ;
  END
END AOI22_X2

MACRO BUF_X1
  CLASS core ;
  FOREIGN BUF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.32 BY 0.768 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.576 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.24 0.114 0.272 0.704 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.1429 0.796 ;
        RECT 0.1429 0.74 0.33 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.33 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.072 0.115 0.185 ;
        RECT 0.114 0.185 0.115 0.213 ;
        RECT 0.114 0.428 0.115 0.456 ;
        RECT 0.114 0.456 0.115 0.558 ;
        RECT 0.115 0.072 0.1419 0.185 ;
        RECT 0.115 0.185 0.1419 0.213 ;
        RECT 0.115 0.213 0.1419 0.428 ;
        RECT 0.115 0.428 0.1419 0.456 ;
        RECT 0.115 0.456 0.1419 0.558 ;
        RECT 0.1419 0.185 0.1429 0.213 ;
        RECT 0.1419 0.213 0.1429 0.428 ;
        RECT 0.1419 0.428 0.1429 0.456 ;
      LAYER M1 ;
        RECT 0.114 0.072 0.115 0.185 ;
        RECT 0.114 0.185 0.115 0.213 ;
        RECT 0.114 0.428 0.115 0.456 ;
        RECT 0.114 0.456 0.115 0.558 ;
        RECT 0.115 0.072 0.1419 0.185 ;
        RECT 0.115 0.185 0.1419 0.213 ;
        RECT 0.115 0.213 0.1419 0.428 ;
        RECT 0.115 0.428 0.1419 0.456 ;
        RECT 0.115 0.456 0.1419 0.558 ;
        RECT 0.1419 0.185 0.1429 0.213 ;
        RECT 0.1419 0.213 0.1429 0.428 ;
        RECT 0.1419 0.428 0.1429 0.456 ;
  END
END BUF_X1

MACRO BUF_X2
  CLASS core ;
  FOREIGN BUF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.32 BY 0.768 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.267 0.078 0.512 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1739 0.603 0.177 0.704 ;
        RECT 0.177 0.072 0.178 0.132 ;
        RECT 0.177 0.603 0.178 0.704 ;
        RECT 0.178 0.072 0.206 0.132 ;
        RECT 0.178 0.132 0.206 0.603 ;
        RECT 0.178 0.603 0.206 0.704 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.1419 0.796 ;
        RECT 0.1419 0.74 0.33 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.33 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.042 0.556 0.05 0.584 ;
        RECT 0.042 0.584 0.05 0.686 ;
        RECT 0.05 0.096 0.078 0.192 ;
        RECT 0.05 0.192 0.078 0.22 ;
        RECT 0.05 0.556 0.078 0.584 ;
        RECT 0.05 0.584 0.078 0.686 ;
        RECT 0.078 0.192 0.0859 0.22 ;
        RECT 0.078 0.556 0.0859 0.584 ;
        RECT 0.078 0.584 0.0859 0.686 ;
        RECT 0.0859 0.192 0.114 0.22 ;
        RECT 0.0859 0.556 0.114 0.584 ;
        RECT 0.114 0.192 0.1419 0.22 ;
        RECT 0.114 0.22 0.1419 0.556 ;
        RECT 0.114 0.556 0.1419 0.584 ;
      LAYER M1 ;
        RECT 0.042 0.556 0.05 0.584 ;
        RECT 0.042 0.584 0.05 0.686 ;
        RECT 0.05 0.096 0.078 0.192 ;
        RECT 0.05 0.192 0.078 0.22 ;
        RECT 0.05 0.556 0.078 0.584 ;
        RECT 0.05 0.584 0.078 0.686 ;
        RECT 0.078 0.192 0.0859 0.22 ;
        RECT 0.078 0.556 0.0859 0.584 ;
        RECT 0.078 0.584 0.0859 0.686 ;
        RECT 0.0859 0.192 0.114 0.22 ;
        RECT 0.0859 0.556 0.114 0.584 ;
        RECT 0.114 0.192 0.1419 0.22 ;
        RECT 0.114 0.22 0.1419 0.556 ;
        RECT 0.114 0.556 0.1419 0.584 ;
  END
END BUF_X2

MACRO BUF_X4
  CLASS core ;
  FOREIGN BUF_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.768 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.242 0.206 0.526 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.145 0.1019 0.21 0.13 ;
        RECT 0.21 0.1019 0.27 0.13 ;
        RECT 0.21 0.638 0.27 0.666 ;
        RECT 0.27 0.1019 0.368 0.13 ;
        RECT 0.27 0.638 0.368 0.666 ;
        RECT 0.368 0.1019 0.4 0.13 ;
        RECT 0.368 0.13 0.4 0.638 ;
        RECT 0.368 0.638 0.4 0.666 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.27 0.796 ;
        RECT 0.27 0.74 0.522 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.522 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.027 0.166 0.0859 0.198 ;
        RECT 0.0859 0.166 0.242 0.198 ;
        RECT 0.0859 0.5699 0.242 0.602 ;
        RECT 0.242 0.166 0.27 0.198 ;
        RECT 0.242 0.198 0.27 0.5699 ;
        RECT 0.242 0.5699 0.27 0.602 ;
      LAYER M1 ;
        RECT 0.027 0.166 0.0859 0.198 ;
        RECT 0.0859 0.166 0.242 0.198 ;
        RECT 0.0859 0.5699 0.242 0.602 ;
        RECT 0.242 0.166 0.27 0.198 ;
        RECT 0.242 0.198 0.27 0.5699 ;
        RECT 0.242 0.5699 0.27 0.602 ;
  END
END BUF_X4

MACRO BUF_X8
  CLASS core ;
  FOREIGN BUF_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.896 BY 0.768 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.366 ;
        RECT 0.05 0.366 0.078 0.398 ;
        RECT 0.05 0.398 0.078 0.512 ;
        RECT 0.078 0.366 0.298 0.398 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.338 0.1019 0.7 0.13 ;
        RECT 0.338 0.638 0.7 0.666 ;
        RECT 0.7 0.1019 0.754 0.13 ;
        RECT 0.7 0.638 0.754 0.666 ;
        RECT 0.754 0.1019 0.782 0.13 ;
        RECT 0.754 0.13 0.782 0.638 ;
        RECT 0.754 0.638 0.782 0.666 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.7 0.796 ;
        RECT 0.7 0.74 0.906 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.906 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.099 0.098 0.114 0.186 ;
        RECT 0.099 0.186 0.114 0.214 ;
        RECT 0.114 0.098 0.1419 0.186 ;
        RECT 0.114 0.186 0.1419 0.214 ;
        RECT 0.114 0.527 0.1419 0.583 ;
        RECT 0.114 0.583 0.1419 0.67 ;
        RECT 0.1419 0.098 0.157 0.186 ;
        RECT 0.1419 0.186 0.157 0.214 ;
        RECT 0.1419 0.527 0.157 0.583 ;
        RECT 0.157 0.186 0.354 0.214 ;
        RECT 0.157 0.527 0.354 0.583 ;
        RECT 0.354 0.186 0.382 0.214 ;
        RECT 0.354 0.214 0.382 0.341 ;
        RECT 0.354 0.341 0.382 0.369 ;
        RECT 0.354 0.369 0.382 0.527 ;
        RECT 0.354 0.527 0.382 0.583 ;
        RECT 0.382 0.341 0.7 0.369 ;
      LAYER M1 ;
        RECT 0.099 0.098 0.114 0.186 ;
        RECT 0.099 0.186 0.114 0.214 ;
        RECT 0.114 0.098 0.1419 0.186 ;
        RECT 0.114 0.186 0.1419 0.214 ;
        RECT 0.114 0.527 0.1419 0.583 ;
        RECT 0.114 0.583 0.1419 0.67 ;
        RECT 0.1419 0.098 0.157 0.186 ;
        RECT 0.1419 0.186 0.157 0.214 ;
        RECT 0.1419 0.527 0.157 0.583 ;
        RECT 0.157 0.186 0.354 0.214 ;
        RECT 0.157 0.527 0.354 0.583 ;
        RECT 0.354 0.186 0.382 0.214 ;
        RECT 0.354 0.214 0.382 0.341 ;
        RECT 0.354 0.341 0.382 0.369 ;
        RECT 0.354 0.369 0.382 0.527 ;
        RECT 0.354 0.527 0.382 0.583 ;
        RECT 0.382 0.341 0.7 0.369 ;
  END
END BUF_X8

MACRO BUF_X12
  CLASS core ;
  FOREIGN BUF_X12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.28 BY 0.768 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.048 0.236 0.08 0.366 ;
        RECT 0.048 0.366 0.08 0.398 ;
        RECT 0.048 0.398 0.08 0.515 ;
        RECT 0.08 0.366 0.426 0.398 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.466 0.1019 1.07 0.13 ;
        RECT 0.466 0.638 1.07 0.666 ;
        RECT 1.07 0.1019 1.1359 0.13 ;
        RECT 1.07 0.638 1.1359 0.666 ;
        RECT 1.1359 0.1019 1.168 0.13 ;
        RECT 1.1359 0.13 1.168 0.638 ;
        RECT 1.1359 0.638 1.168 0.666 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.07 0.796 ;
        RECT 1.07 0.74 1.29 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.29 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.098 0.551 0.112 0.583 ;
        RECT 0.098 0.583 0.112 0.67 ;
        RECT 0.112 0.098 0.144 0.185 ;
        RECT 0.112 0.185 0.144 0.217 ;
        RECT 0.112 0.551 0.144 0.583 ;
        RECT 0.112 0.583 0.144 0.67 ;
        RECT 0.144 0.185 0.157 0.217 ;
        RECT 0.144 0.551 0.157 0.583 ;
        RECT 0.144 0.583 0.157 0.67 ;
        RECT 0.157 0.185 0.462 0.217 ;
        RECT 0.157 0.551 0.462 0.583 ;
        RECT 0.462 0.185 0.49 0.217 ;
        RECT 0.462 0.217 0.49 0.37 ;
        RECT 0.462 0.37 0.49 0.398 ;
        RECT 0.462 0.398 0.49 0.551 ;
        RECT 0.462 0.551 0.49 0.583 ;
        RECT 0.49 0.37 1.07 0.398 ;
      LAYER M1 ;
        RECT 0.098 0.551 0.112 0.583 ;
        RECT 0.098 0.583 0.112 0.67 ;
        RECT 0.112 0.098 0.144 0.185 ;
        RECT 0.112 0.185 0.144 0.217 ;
        RECT 0.112 0.551 0.144 0.583 ;
        RECT 0.112 0.583 0.144 0.67 ;
        RECT 0.144 0.185 0.157 0.217 ;
        RECT 0.144 0.551 0.157 0.583 ;
        RECT 0.144 0.583 0.157 0.67 ;
        RECT 0.157 0.185 0.462 0.217 ;
        RECT 0.157 0.551 0.462 0.583 ;
        RECT 0.462 0.185 0.49 0.217 ;
        RECT 0.462 0.217 0.49 0.37 ;
        RECT 0.462 0.37 0.49 0.398 ;
        RECT 0.462 0.398 0.49 0.551 ;
        RECT 0.462 0.551 0.49 0.583 ;
        RECT 0.49 0.37 1.07 0.398 ;
  END
END BUF_X12

MACRO BUF_X16
  CLASS core ;
  FOREIGN BUF_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.664 BY 0.768 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.232 0.078 0.355 ;
        RECT 0.05 0.355 0.078 0.413 ;
        RECT 0.05 0.413 0.078 0.512 ;
        RECT 0.078 0.355 0.554 0.413 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.594 0.1019 1.454 0.13 ;
        RECT 0.594 0.632 1.454 0.66 ;
        RECT 1.454 0.1019 1.52 0.13 ;
        RECT 1.454 0.632 1.52 0.66 ;
        RECT 1.52 0.1019 1.552 0.13 ;
        RECT 1.52 0.13 1.552 0.632 ;
        RECT 1.52 0.632 1.552 0.66 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.454 0.796 ;
        RECT 1.454 0.74 1.674 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.674 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.098 0.1419 0.205 ;
        RECT 0.114 0.205 0.1419 0.233 ;
        RECT 0.114 0.458 0.1419 0.486 ;
        RECT 0.114 0.486 0.1419 0.643 ;
        RECT 0.1419 0.205 0.59 0.233 ;
        RECT 0.1419 0.458 0.59 0.486 ;
        RECT 0.59 0.205 0.618 0.233 ;
        RECT 0.59 0.233 0.618 0.368 ;
        RECT 0.59 0.368 0.618 0.396 ;
        RECT 0.59 0.396 0.618 0.458 ;
        RECT 0.59 0.458 0.618 0.486 ;
        RECT 0.618 0.368 1.454 0.396 ;
      LAYER M1 ;
        RECT 0.114 0.098 0.1419 0.205 ;
        RECT 0.114 0.205 0.1419 0.233 ;
        RECT 0.114 0.458 0.1419 0.486 ;
        RECT 0.114 0.486 0.1419 0.643 ;
        RECT 0.1419 0.205 0.59 0.233 ;
        RECT 0.1419 0.458 0.59 0.486 ;
        RECT 0.59 0.205 0.618 0.233 ;
        RECT 0.59 0.233 0.618 0.368 ;
        RECT 0.59 0.368 0.618 0.396 ;
        RECT 0.59 0.396 0.618 0.458 ;
        RECT 0.59 0.458 0.618 0.486 ;
        RECT 0.618 0.368 1.454 0.396 ;
  END
END BUF_X16

MACRO CLKBUF_X1
  CLASS core ;
  FOREIGN CLKBUF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.32 BY 0.768 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.576 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.24 0.114 0.272 0.704 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.1429 0.796 ;
        RECT 0.1429 0.74 0.33 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.33 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.072 0.115 0.185 ;
        RECT 0.114 0.185 0.115 0.213 ;
        RECT 0.114 0.393 0.115 0.458 ;
        RECT 0.114 0.458 0.115 0.523 ;
        RECT 0.115 0.072 0.1419 0.185 ;
        RECT 0.115 0.185 0.1419 0.213 ;
        RECT 0.115 0.213 0.1419 0.393 ;
        RECT 0.115 0.393 0.1419 0.458 ;
        RECT 0.115 0.458 0.1419 0.523 ;
        RECT 0.1419 0.185 0.1429 0.213 ;
        RECT 0.1419 0.213 0.1429 0.393 ;
        RECT 0.1419 0.393 0.1429 0.458 ;
      LAYER M1 ;
        RECT 0.114 0.072 0.115 0.185 ;
        RECT 0.114 0.185 0.115 0.213 ;
        RECT 0.114 0.393 0.115 0.458 ;
        RECT 0.114 0.458 0.115 0.523 ;
        RECT 0.115 0.072 0.1419 0.185 ;
        RECT 0.115 0.185 0.1419 0.213 ;
        RECT 0.115 0.213 0.1419 0.393 ;
        RECT 0.115 0.393 0.1419 0.458 ;
        RECT 0.115 0.458 0.1419 0.523 ;
        RECT 0.1419 0.185 0.1429 0.213 ;
        RECT 0.1419 0.213 0.1429 0.393 ;
        RECT 0.1419 0.393 0.1429 0.458 ;
  END
END CLKBUF_X1

MACRO CLKBUF_X2
  CLASS core ;
  FOREIGN CLKBUF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.32 BY 0.768 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.296 0.078 0.512 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1739 0.638 0.178 0.704 ;
        RECT 0.178 0.072 0.206 0.638 ;
        RECT 0.178 0.638 0.206 0.704 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.1419 0.796 ;
        RECT 0.1419 0.74 0.33 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.33 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.129 0.08 0.192 ;
        RECT 0.048 0.192 0.08 0.22 ;
        RECT 0.048 0.556 0.08 0.584 ;
        RECT 0.048 0.584 0.08 0.686 ;
        RECT 0.08 0.192 0.114 0.22 ;
        RECT 0.08 0.556 0.114 0.584 ;
        RECT 0.114 0.192 0.1419 0.22 ;
        RECT 0.114 0.22 0.1419 0.556 ;
        RECT 0.114 0.556 0.1419 0.584 ;
      LAYER M1 ;
        RECT 0.048 0.129 0.08 0.192 ;
        RECT 0.048 0.192 0.08 0.22 ;
        RECT 0.048 0.556 0.08 0.584 ;
        RECT 0.048 0.584 0.08 0.686 ;
        RECT 0.08 0.192 0.114 0.22 ;
        RECT 0.08 0.556 0.114 0.584 ;
        RECT 0.114 0.192 0.1419 0.22 ;
        RECT 0.114 0.22 0.1419 0.556 ;
        RECT 0.114 0.556 0.1419 0.584 ;
  END
END CLKBUF_X2

MACRO CLKBUF_X4
  CLASS core ;
  FOREIGN CLKBUF_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.768 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.242 0.1419 0.526 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.145 0.1019 0.205 0.13 ;
        RECT 0.205 0.1019 0.206 0.13 ;
        RECT 0.205 0.638 0.206 0.666 ;
        RECT 0.206 0.1019 0.368 0.13 ;
        RECT 0.206 0.638 0.368 0.666 ;
        RECT 0.368 0.1019 0.4 0.13 ;
        RECT 0.368 0.13 0.4 0.638 ;
        RECT 0.368 0.638 0.4 0.666 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.206 0.796 ;
        RECT 0.206 0.74 0.522 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.522 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.041 0.166 0.082 0.194 ;
        RECT 0.082 0.166 0.178 0.194 ;
        RECT 0.082 0.574 0.178 0.602 ;
        RECT 0.178 0.166 0.206 0.194 ;
        RECT 0.178 0.194 0.206 0.574 ;
        RECT 0.178 0.574 0.206 0.602 ;
      LAYER M1 ;
        RECT 0.041 0.166 0.082 0.194 ;
        RECT 0.082 0.166 0.178 0.194 ;
        RECT 0.082 0.574 0.178 0.602 ;
        RECT 0.178 0.166 0.206 0.194 ;
        RECT 0.178 0.194 0.206 0.574 ;
        RECT 0.178 0.574 0.206 0.602 ;
  END
END CLKBUF_X4

MACRO CLKBUF_X8
  CLASS core ;
  FOREIGN CLKBUF_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.896 BY 0.768 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.328 ;
        RECT 0.05 0.328 0.078 0.356 ;
        RECT 0.05 0.356 0.078 0.512 ;
        RECT 0.078 0.256 0.079 0.328 ;
        RECT 0.078 0.328 0.079 0.356 ;
        RECT 0.079 0.328 0.318 0.356 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.338 0.1019 0.718 0.13 ;
        RECT 0.338 0.638 0.718 0.666 ;
        RECT 0.718 0.1019 0.754 0.13 ;
        RECT 0.718 0.638 0.754 0.666 ;
        RECT 0.754 0.1019 0.782 0.13 ;
        RECT 0.754 0.13 0.782 0.638 ;
        RECT 0.754 0.638 0.782 0.666 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.718 0.796 ;
        RECT 0.718 0.74 0.906 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.906 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.166 0.114 0.194 ;
        RECT 0.114 0.166 0.1419 0.194 ;
        RECT 0.114 0.45 0.1419 0.482 ;
        RECT 0.114 0.482 0.1419 0.542 ;
        RECT 0.1419 0.166 0.406 0.194 ;
        RECT 0.1419 0.45 0.406 0.482 ;
        RECT 0.406 0.166 0.434 0.194 ;
        RECT 0.406 0.194 0.434 0.357 ;
        RECT 0.406 0.357 0.434 0.415 ;
        RECT 0.406 0.415 0.434 0.45 ;
        RECT 0.406 0.45 0.434 0.482 ;
        RECT 0.434 0.357 0.718 0.415 ;
      LAYER M1 ;
        RECT 0.05 0.166 0.114 0.194 ;
        RECT 0.114 0.166 0.1419 0.194 ;
        RECT 0.114 0.45 0.1419 0.482 ;
        RECT 0.114 0.482 0.1419 0.542 ;
        RECT 0.1419 0.166 0.406 0.194 ;
        RECT 0.1419 0.45 0.406 0.482 ;
        RECT 0.406 0.166 0.434 0.194 ;
        RECT 0.406 0.194 0.434 0.357 ;
        RECT 0.406 0.357 0.434 0.415 ;
        RECT 0.406 0.415 0.434 0.45 ;
        RECT 0.406 0.45 0.434 0.482 ;
        RECT 0.434 0.357 0.718 0.415 ;
  END
END CLKBUF_X8

MACRO CLKBUF_X12
  CLASS core ;
  FOREIGN CLKBUF_X12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.28 BY 0.768 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.238 0.083 0.336 ;
        RECT 0.045 0.336 0.083 0.368 ;
        RECT 0.045 0.368 0.083 0.53 ;
        RECT 0.083 0.336 0.426 0.368 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.466 0.1019 0.998 0.13 ;
        RECT 0.466 0.638 0.998 0.666 ;
        RECT 0.998 0.1019 1.1359 0.13 ;
        RECT 0.998 0.638 1.1359 0.666 ;
        RECT 1.1359 0.1019 1.168 0.13 ;
        RECT 1.1359 0.13 1.168 0.638 ;
        RECT 1.1359 0.638 1.168 0.666 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.998 0.796 ;
        RECT 0.998 0.74 1.29 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.29 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.0429 0.166 0.114 0.194 ;
        RECT 0.114 0.166 0.1419 0.194 ;
        RECT 0.114 0.55 0.1419 0.578 ;
        RECT 0.114 0.578 0.1419 0.67 ;
        RECT 0.1419 0.166 0.462 0.194 ;
        RECT 0.1419 0.55 0.462 0.578 ;
        RECT 0.462 0.166 0.49 0.194 ;
        RECT 0.462 0.194 0.49 0.314 ;
        RECT 0.462 0.314 0.49 0.3459 ;
        RECT 0.462 0.3459 0.49 0.55 ;
        RECT 0.462 0.55 0.49 0.578 ;
        RECT 0.49 0.166 0.494 0.194 ;
        RECT 0.49 0.194 0.494 0.314 ;
        RECT 0.49 0.314 0.494 0.3459 ;
        RECT 0.494 0.314 0.998 0.3459 ;
      LAYER M1 ;
        RECT 0.0429 0.166 0.114 0.194 ;
        RECT 0.114 0.166 0.1419 0.194 ;
        RECT 0.114 0.55 0.1419 0.578 ;
        RECT 0.114 0.578 0.1419 0.67 ;
        RECT 0.1419 0.166 0.462 0.194 ;
        RECT 0.1419 0.55 0.462 0.578 ;
        RECT 0.462 0.166 0.49 0.194 ;
        RECT 0.462 0.194 0.49 0.314 ;
        RECT 0.462 0.314 0.49 0.3459 ;
        RECT 0.462 0.3459 0.49 0.55 ;
        RECT 0.462 0.55 0.49 0.578 ;
        RECT 0.49 0.166 0.494 0.194 ;
        RECT 0.49 0.194 0.494 0.314 ;
        RECT 0.49 0.314 0.494 0.3459 ;
        RECT 0.494 0.314 0.998 0.3459 ;
  END
END CLKBUF_X12

MACRO CLKBUF_X16
  CLASS core ;
  FOREIGN CLKBUF_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.664 BY 0.768 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.222 0.078 0.326 ;
        RECT 0.05 0.326 0.078 0.358 ;
        RECT 0.05 0.358 0.078 0.526 ;
        RECT 0.078 0.326 0.554 0.358 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.594 0.0869 1.454 0.145 ;
        RECT 0.594 0.623 1.454 0.681 ;
        RECT 1.454 0.0869 1.52 0.145 ;
        RECT 1.454 0.623 1.52 0.681 ;
        RECT 1.52 0.0869 1.552 0.145 ;
        RECT 1.52 0.145 1.552 0.623 ;
        RECT 1.52 0.623 1.552 0.681 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.454 0.796 ;
        RECT 1.454 0.74 1.674 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.674 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.109 0.1419 0.205 ;
        RECT 0.114 0.205 0.1419 0.233 ;
        RECT 0.114 0.525 0.1419 0.5629 ;
        RECT 0.114 0.5629 0.1419 0.638 ;
        RECT 0.1419 0.205 0.595 0.233 ;
        RECT 0.1419 0.525 0.595 0.5629 ;
        RECT 0.595 0.205 0.653 0.233 ;
        RECT 0.595 0.233 0.653 0.316 ;
        RECT 0.595 0.316 0.653 0.3439 ;
        RECT 0.595 0.3439 0.653 0.525 ;
        RECT 0.595 0.525 0.653 0.5629 ;
        RECT 0.653 0.316 1.454 0.3439 ;
      LAYER M1 ;
        RECT 0.114 0.109 0.1419 0.205 ;
        RECT 0.114 0.205 0.1419 0.233 ;
        RECT 0.114 0.525 0.1419 0.5629 ;
        RECT 0.114 0.5629 0.1419 0.638 ;
        RECT 0.1419 0.205 0.595 0.233 ;
        RECT 0.1419 0.525 0.595 0.5629 ;
        RECT 0.595 0.205 0.653 0.233 ;
        RECT 0.595 0.233 0.653 0.316 ;
        RECT 0.595 0.316 0.653 0.3439 ;
        RECT 0.595 0.3439 0.653 0.525 ;
        RECT 0.595 0.525 0.653 0.5629 ;
        RECT 0.653 0.316 1.454 0.3439 ;
  END
END CLKBUF_X16

MACRO CLKGATETST_X1
  CLASS core ;
  FOREIGN CLKGATETST_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.088 BY 0.768 ;
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.6899 0.238 0.718 0.512 ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.1419 0.672 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.32 0.078 0.672 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.01 0.096 1.038 0.654 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.366 0.796 ;
        RECT 0.366 0.74 0.91 0.796 ;
        RECT 0.91 0.74 0.974 0.796 ;
        RECT 0.974 0.74 1.098 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.098 0.028 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.21 0.402 0.686 0.43 ;
        RECT 0.146 0.466 0.522 0.494 ;
        RECT 0.73 0.402 1.006 0.43 ;
      LAYER MINT1 ;
        RECT 0.21 0.402 0.686 0.43 ;
        RECT 0.146 0.466 0.522 0.494 ;
        RECT 0.73 0.402 1.006 0.43 ;
      LAYER M1 ;
        RECT 0.048 0.1019 0.08 0.13 ;
        RECT 0.048 0.13 0.08 0.213 ;
        RECT 0.08 0.1019 0.238 0.13 ;
        RECT 0.242 0.264 0.27 0.541 ;
        RECT 0.37 0.242 0.398 0.502 ;
        RECT 0.462 0.372 0.494 0.51 ;
        RECT 0.626 0.166 0.654 0.194 ;
        RECT 0.626 0.194 0.654 0.556 ;
        RECT 0.626 0.556 0.654 0.592 ;
        RECT 0.654 0.166 0.75 0.194 ;
        RECT 0.654 0.556 0.75 0.592 ;
        RECT 0.75 0.166 0.755 0.194 ;
        RECT 0.754 0.248 0.79 0.463 ;
        RECT 0.754 0.463 0.79 0.502 ;
        RECT 0.79 0.463 0.8179 0.502 ;
        RECT 0.8179 0.463 0.846 0.502 ;
        RECT 0.8179 0.502 0.846 0.584 ;
        RECT 0.946 0.226 0.974 0.574 ;
        RECT 0.178 0.166 0.206 0.194 ;
        RECT 0.178 0.194 0.206 0.628 ;
        RECT 0.178 0.628 0.206 0.676 ;
        RECT 0.206 0.166 0.302 0.194 ;
        RECT 0.206 0.628 0.302 0.676 ;
        RECT 0.302 0.628 0.366 0.676 ;
        RECT 0.306 0.307 0.334 0.546 ;
        RECT 0.306 0.546 0.334 0.574 ;
        RECT 0.334 0.546 0.558 0.574 ;
        RECT 0.558 0.184 0.59 0.307 ;
        RECT 0.558 0.307 0.59 0.546 ;
        RECT 0.558 0.546 0.59 0.574 ;
        RECT 0.434 0.1019 0.462 0.13 ;
        RECT 0.434 0.13 0.462 0.334 ;
        RECT 0.462 0.1019 0.466 0.13 ;
        RECT 0.466 0.1019 0.882 0.13 ;
        RECT 0.466 0.628 0.882 0.676 ;
        RECT 0.882 0.1019 0.91 0.13 ;
        RECT 0.882 0.13 0.91 0.334 ;
        RECT 0.882 0.334 0.91 0.628 ;
        RECT 0.882 0.628 0.91 0.676 ;
      LAYER V1 ;
        RECT 0.178 0.466 0.206 0.494 ;
        RECT 0.242 0.402 0.27 0.43 ;
        RECT 0.37 0.402 0.398 0.43 ;
        RECT 0.462 0.466 0.49 0.494 ;
        RECT 0.626 0.402 0.654 0.43 ;
        RECT 0.762 0.402 0.79 0.43 ;
        RECT 0.946 0.402 0.974 0.43 ;
      LAYER M1 ;
        RECT 0.048 0.1019 0.08 0.13 ;
        RECT 0.048 0.13 0.08 0.213 ;
        RECT 0.08 0.1019 0.238 0.13 ;
        RECT 0.242 0.264 0.27 0.541 ;
        RECT 0.37 0.242 0.398 0.502 ;
        RECT 0.462 0.372 0.494 0.51 ;
        RECT 0.626 0.166 0.654 0.194 ;
        RECT 0.626 0.194 0.654 0.556 ;
        RECT 0.626 0.556 0.654 0.592 ;
        RECT 0.654 0.166 0.75 0.194 ;
        RECT 0.654 0.556 0.75 0.592 ;
        RECT 0.75 0.166 0.755 0.194 ;
        RECT 0.754 0.248 0.79 0.463 ;
        RECT 0.754 0.463 0.79 0.502 ;
        RECT 0.79 0.463 0.8179 0.502 ;
        RECT 0.8179 0.463 0.846 0.502 ;
        RECT 0.8179 0.502 0.846 0.584 ;
        RECT 0.946 0.226 0.974 0.574 ;
        RECT 0.178 0.166 0.206 0.194 ;
        RECT 0.178 0.194 0.206 0.628 ;
        RECT 0.178 0.628 0.206 0.676 ;
        RECT 0.206 0.166 0.302 0.194 ;
        RECT 0.206 0.628 0.302 0.676 ;
        RECT 0.302 0.628 0.366 0.676 ;
        RECT 0.306 0.307 0.334 0.546 ;
        RECT 0.306 0.546 0.334 0.574 ;
        RECT 0.334 0.546 0.558 0.574 ;
        RECT 0.558 0.184 0.59 0.307 ;
        RECT 0.558 0.307 0.59 0.546 ;
        RECT 0.558 0.546 0.59 0.574 ;
        RECT 0.434 0.1019 0.462 0.13 ;
        RECT 0.434 0.13 0.462 0.334 ;
        RECT 0.462 0.1019 0.466 0.13 ;
        RECT 0.466 0.1019 0.882 0.13 ;
        RECT 0.466 0.628 0.882 0.676 ;
        RECT 0.882 0.1019 0.91 0.13 ;
        RECT 0.882 0.13 0.91 0.334 ;
        RECT 0.882 0.334 0.91 0.628 ;
        RECT 0.882 0.628 0.91 0.676 ;
  END
END CLKGATETST_X1

MACRO DFFRNQ_X1
  CLASS core ;
  FOREIGN DFFRNQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.664 BY 0.768 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.242 0.27 0.526 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.704 0.274 1.1339 0.302 ;
        RECT 1.1339 0.274 1.326 0.302 ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.512 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.064 1.616 0.704 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.1419 0.796 ;
        RECT 0.1419 0.74 0.206 0.796 ;
        RECT 0.206 0.74 0.334 0.796 ;
        RECT 0.334 0.74 0.398 0.796 ;
        RECT 0.398 0.74 0.526 0.796 ;
        RECT 0.526 0.74 0.8139 0.796 ;
        RECT 0.8139 0.74 0.91 0.796 ;
        RECT 0.91 0.74 0.974 0.796 ;
        RECT 0.974 0.74 1.102 0.796 ;
        RECT 1.102 0.74 1.188 0.796 ;
        RECT 1.188 0.74 1.488 0.796 ;
        RECT 1.488 0.74 1.674 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.674 0.028 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.146 0.21 1.1339 0.238 ;
        RECT 0.082 0.53 1.1339 0.558 ;
      LAYER MINT1 ;
        RECT 0.146 0.21 1.1339 0.238 ;
        RECT 0.082 0.53 1.1339 0.558 ;
      LAYER M1 ;
        RECT 0.178 0.072 0.206 0.6959 ;
        RECT 0.306 0.072 0.334 0.6959 ;
        RECT 0.53 0.623 0.8139 0.681 ;
        RECT 0.434 0.1019 0.462 0.13 ;
        RECT 0.434 0.13 0.462 0.438 ;
        RECT 0.434 0.438 0.462 0.67 ;
        RECT 0.462 0.1019 0.8 0.13 ;
        RECT 0.8 0.1019 0.828 0.13 ;
        RECT 0.8 0.13 0.828 0.438 ;
        RECT 0.576 0.33 0.604 0.506 ;
        RECT 0.576 0.506 0.604 0.534 ;
        RECT 0.604 0.506 0.882 0.534 ;
        RECT 0.882 0.072 0.91 0.33 ;
        RECT 0.882 0.33 0.91 0.506 ;
        RECT 0.882 0.506 0.91 0.534 ;
        RECT 0.882 0.534 0.91 0.672 ;
        RECT 1.01 0.1019 1.038 0.13 ;
        RECT 1.01 0.13 1.038 0.366 ;
        RECT 1.01 0.366 1.038 0.67 ;
        RECT 1.038 0.1019 1.335 0.13 ;
        RECT 1.335 0.1019 1.363 0.13 ;
        RECT 1.335 0.13 1.363 0.366 ;
        RECT 1.224 0.394 1.252 0.638 ;
        RECT 1.224 0.638 1.252 0.666 ;
        RECT 1.252 0.638 1.458 0.666 ;
        RECT 1.458 0.072 1.486 0.132 ;
        RECT 1.458 0.132 1.486 0.394 ;
        RECT 1.458 0.394 1.486 0.638 ;
        RECT 1.458 0.638 1.486 0.666 ;
        RECT 1.486 0.132 1.488 0.394 ;
        RECT 1.486 0.394 1.488 0.638 ;
        RECT 1.486 0.638 1.488 0.666 ;
        RECT 0.048 0.085 0.08 0.1409 ;
        RECT 0.048 0.1409 0.08 0.169 ;
        RECT 0.048 0.5669 0.08 0.606 ;
        RECT 0.048 0.606 0.08 0.686 ;
        RECT 0.08 0.1409 0.114 0.169 ;
        RECT 0.08 0.5669 0.114 0.606 ;
        RECT 0.114 0.1409 0.1419 0.169 ;
        RECT 0.114 0.169 0.1419 0.5669 ;
        RECT 0.114 0.5669 0.1419 0.606 ;
        RECT 0.37 0.194 0.398 0.494 ;
        RECT 0.498 0.402 0.526 0.574 ;
        RECT 0.526 0.194 0.558 0.294 ;
        RECT 0.736 0.258 0.764 0.438 ;
        RECT 0.946 0.274 0.974 0.578 ;
        RECT 1.074 0.1739 1.102 0.317 ;
        RECT 1.074 0.46 1.102 0.622 ;
        RECT 1.156 0.166 1.188 0.686 ;
        RECT 1.266 0.1739 1.294 0.318 ;
      LAYER V1 ;
        RECT 0.114 0.53 0.1419 0.558 ;
        RECT 0.178 0.21 0.206 0.238 ;
        RECT 0.37 0.21 0.398 0.238 ;
        RECT 0.498 0.53 0.526 0.558 ;
        RECT 0.53 0.21 0.558 0.238 ;
        RECT 0.736 0.274 0.764 0.302 ;
        RECT 0.946 0.53 0.974 0.558 ;
        RECT 1.074 0.21 1.102 0.238 ;
        RECT 1.074 0.53 1.102 0.558 ;
        RECT 1.266 0.274 1.294 0.302 ;
      LAYER M1 ;
        RECT 0.178 0.072 0.206 0.6959 ;
        RECT 0.306 0.072 0.334 0.6959 ;
        RECT 0.53 0.623 0.8139 0.681 ;
        RECT 0.434 0.1019 0.462 0.13 ;
        RECT 0.434 0.13 0.462 0.438 ;
        RECT 0.434 0.438 0.462 0.67 ;
        RECT 0.462 0.1019 0.8 0.13 ;
        RECT 0.8 0.1019 0.828 0.13 ;
        RECT 0.8 0.13 0.828 0.438 ;
        RECT 0.576 0.33 0.604 0.506 ;
        RECT 0.576 0.506 0.604 0.534 ;
        RECT 0.604 0.506 0.882 0.534 ;
        RECT 0.882 0.072 0.91 0.33 ;
        RECT 0.882 0.33 0.91 0.506 ;
        RECT 0.882 0.506 0.91 0.534 ;
        RECT 0.882 0.534 0.91 0.672 ;
        RECT 1.01 0.1019 1.038 0.13 ;
        RECT 1.01 0.13 1.038 0.366 ;
        RECT 1.01 0.366 1.038 0.67 ;
        RECT 1.038 0.1019 1.335 0.13 ;
        RECT 1.335 0.1019 1.363 0.13 ;
        RECT 1.335 0.13 1.363 0.366 ;
        RECT 1.224 0.394 1.252 0.638 ;
        RECT 1.224 0.638 1.252 0.666 ;
        RECT 1.252 0.638 1.458 0.666 ;
        RECT 1.458 0.072 1.486 0.132 ;
        RECT 1.458 0.132 1.486 0.394 ;
        RECT 1.458 0.394 1.486 0.638 ;
        RECT 1.458 0.638 1.486 0.666 ;
        RECT 1.486 0.132 1.488 0.394 ;
        RECT 1.486 0.394 1.488 0.638 ;
        RECT 1.486 0.638 1.488 0.666 ;
        RECT 0.048 0.085 0.08 0.1409 ;
        RECT 0.048 0.1409 0.08 0.169 ;
        RECT 0.048 0.5669 0.08 0.606 ;
        RECT 0.048 0.606 0.08 0.686 ;
        RECT 0.08 0.1409 0.114 0.169 ;
        RECT 0.08 0.5669 0.114 0.606 ;
        RECT 0.114 0.1409 0.1419 0.169 ;
        RECT 0.114 0.169 0.1419 0.5669 ;
        RECT 0.114 0.5669 0.1419 0.606 ;
        RECT 0.37 0.194 0.398 0.494 ;
        RECT 0.498 0.402 0.526 0.574 ;
        RECT 0.526 0.194 0.558 0.294 ;
        RECT 0.736 0.258 0.764 0.438 ;
        RECT 0.946 0.274 0.974 0.578 ;
        RECT 1.074 0.1739 1.102 0.317 ;
        RECT 1.074 0.46 1.102 0.622 ;
        RECT 1.156 0.166 1.188 0.686 ;
        RECT 1.266 0.1739 1.294 0.318 ;
  END
END DFFRNQ_X1

MACRO DFFSNQ_X1
  CLASS core ;
  FOREIGN DFFSNQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.664 BY 0.768 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.242 0.27 0.526 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.722 0.274 1.1339 0.302 ;
        RECT 1.1339 0.274 1.326 0.302 ;
    END
  END SN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.512 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.064 1.616 0.704 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.1419 0.796 ;
        RECT 0.1419 0.74 0.206 0.796 ;
        RECT 0.206 0.74 0.334 0.796 ;
        RECT 0.334 0.74 0.398 0.796 ;
        RECT 0.398 0.74 0.526 0.796 ;
        RECT 0.526 0.74 0.554 0.796 ;
        RECT 0.554 0.74 0.91 0.796 ;
        RECT 0.91 0.74 0.974 0.796 ;
        RECT 0.974 0.74 1.106 0.796 ;
        RECT 1.106 0.74 1.3899 0.796 ;
        RECT 1.3899 0.74 1.488 0.796 ;
        RECT 1.488 0.74 1.674 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.674 0.028 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.146 0.21 1.1339 0.238 ;
        RECT 0.082 0.53 1.1339 0.558 ;
      LAYER MINT1 ;
        RECT 0.146 0.21 1.1339 0.238 ;
        RECT 0.082 0.53 1.1339 0.558 ;
      LAYER M1 ;
        RECT 0.178 0.072 0.206 0.6959 ;
        RECT 0.306 0.072 0.334 0.6959 ;
        RECT 0.434 0.122 0.462 0.15 ;
        RECT 0.434 0.15 0.462 0.366 ;
        RECT 0.434 0.366 0.462 0.67 ;
        RECT 0.462 0.122 0.8179 0.15 ;
        RECT 0.8179 0.122 0.846 0.15 ;
        RECT 0.8179 0.15 0.846 0.366 ;
        RECT 0.946 0.274 0.974 0.574 ;
        RECT 1.074 0.194 1.106 0.325 ;
        RECT 1.074 0.393 1.106 0.594 ;
        RECT 1.266 0.186 1.294 0.318 ;
        RECT 1.202 0.394 1.23 0.574 ;
        RECT 1.202 0.574 1.23 0.602 ;
        RECT 1.23 0.574 1.458 0.602 ;
        RECT 1.458 0.072 1.486 0.132 ;
        RECT 1.458 0.132 1.486 0.394 ;
        RECT 1.458 0.394 1.486 0.574 ;
        RECT 1.458 0.574 1.486 0.602 ;
        RECT 1.486 0.132 1.488 0.394 ;
        RECT 1.486 0.394 1.488 0.574 ;
        RECT 1.486 0.574 1.488 0.602 ;
        RECT 0.045 0.082 0.048 0.138 ;
        RECT 0.045 0.138 0.048 0.177 ;
        RECT 0.048 0.082 0.08 0.138 ;
        RECT 0.048 0.138 0.08 0.177 ;
        RECT 0.048 0.5669 0.08 0.606 ;
        RECT 0.048 0.606 0.08 0.686 ;
        RECT 0.08 0.082 0.083 0.138 ;
        RECT 0.08 0.138 0.083 0.177 ;
        RECT 0.08 0.5669 0.083 0.606 ;
        RECT 0.083 0.138 0.114 0.177 ;
        RECT 0.083 0.5669 0.114 0.606 ;
        RECT 0.114 0.138 0.1419 0.177 ;
        RECT 0.114 0.177 0.1419 0.5669 ;
        RECT 0.114 0.5669 0.1419 0.606 ;
        RECT 0.37 0.194 0.398 0.494 ;
        RECT 0.498 0.402 0.526 0.59 ;
        RECT 0.526 0.194 0.554 0.305 ;
        RECT 0.754 0.258 0.782 0.366 ;
        RECT 0.608 0.274 0.636 0.574 ;
        RECT 0.608 0.574 0.636 0.602 ;
        RECT 0.636 0.574 0.878 0.602 ;
        RECT 0.878 0.574 0.882 0.602 ;
        RECT 0.878 0.602 0.882 0.686 ;
        RECT 0.882 0.096 0.91 0.274 ;
        RECT 0.882 0.274 0.91 0.574 ;
        RECT 0.882 0.574 0.91 0.602 ;
        RECT 0.882 0.602 0.91 0.686 ;
        RECT 1.01 0.114 1.038 0.1419 ;
        RECT 1.01 0.1419 1.038 0.366 ;
        RECT 1.01 0.366 1.038 0.672 ;
        RECT 1.038 0.114 1.352 0.1419 ;
        RECT 1.352 0.114 1.3799 0.1419 ;
        RECT 1.352 0.1419 1.3799 0.366 ;
        RECT 1.106 0.638 1.3899 0.666 ;
      LAYER V1 ;
        RECT 0.114 0.53 0.1419 0.558 ;
        RECT 0.178 0.21 0.206 0.238 ;
        RECT 0.37 0.21 0.398 0.238 ;
        RECT 0.498 0.53 0.526 0.558 ;
        RECT 0.526 0.21 0.554 0.238 ;
        RECT 0.754 0.274 0.782 0.302 ;
        RECT 0.946 0.53 0.974 0.558 ;
        RECT 1.074 0.21 1.102 0.238 ;
        RECT 1.074 0.53 1.102 0.558 ;
        RECT 1.266 0.274 1.294 0.302 ;
      LAYER M1 ;
        RECT 0.178 0.072 0.206 0.6959 ;
        RECT 0.306 0.072 0.334 0.6959 ;
        RECT 0.434 0.122 0.462 0.15 ;
        RECT 0.434 0.15 0.462 0.366 ;
        RECT 0.434 0.366 0.462 0.67 ;
        RECT 0.462 0.122 0.8179 0.15 ;
        RECT 0.8179 0.122 0.846 0.15 ;
        RECT 0.8179 0.15 0.846 0.366 ;
        RECT 0.946 0.274 0.974 0.574 ;
        RECT 1.074 0.194 1.106 0.325 ;
        RECT 1.074 0.393 1.106 0.594 ;
        RECT 1.266 0.186 1.294 0.318 ;
        RECT 1.202 0.394 1.23 0.574 ;
        RECT 1.202 0.574 1.23 0.602 ;
        RECT 1.23 0.574 1.458 0.602 ;
        RECT 1.458 0.072 1.486 0.132 ;
        RECT 1.458 0.132 1.486 0.394 ;
        RECT 1.458 0.394 1.486 0.574 ;
        RECT 1.458 0.574 1.486 0.602 ;
        RECT 1.486 0.132 1.488 0.394 ;
        RECT 1.486 0.394 1.488 0.574 ;
        RECT 1.486 0.574 1.488 0.602 ;
        RECT 0.045 0.082 0.048 0.138 ;
        RECT 0.045 0.138 0.048 0.177 ;
        RECT 0.048 0.082 0.08 0.138 ;
        RECT 0.048 0.138 0.08 0.177 ;
        RECT 0.048 0.5669 0.08 0.606 ;
        RECT 0.048 0.606 0.08 0.686 ;
        RECT 0.08 0.082 0.083 0.138 ;
        RECT 0.08 0.138 0.083 0.177 ;
        RECT 0.08 0.5669 0.083 0.606 ;
        RECT 0.083 0.138 0.114 0.177 ;
        RECT 0.083 0.5669 0.114 0.606 ;
        RECT 0.114 0.138 0.1419 0.177 ;
        RECT 0.114 0.177 0.1419 0.5669 ;
        RECT 0.114 0.5669 0.1419 0.606 ;
        RECT 0.37 0.194 0.398 0.494 ;
        RECT 0.498 0.402 0.526 0.59 ;
        RECT 0.526 0.194 0.554 0.305 ;
        RECT 0.754 0.258 0.782 0.366 ;
        RECT 0.608 0.274 0.636 0.574 ;
        RECT 0.608 0.574 0.636 0.602 ;
        RECT 0.636 0.574 0.878 0.602 ;
        RECT 0.878 0.574 0.882 0.602 ;
        RECT 0.878 0.602 0.882 0.686 ;
        RECT 0.882 0.096 0.91 0.274 ;
        RECT 0.882 0.274 0.91 0.574 ;
        RECT 0.882 0.574 0.91 0.602 ;
        RECT 0.882 0.602 0.91 0.686 ;
        RECT 1.01 0.114 1.038 0.1419 ;
        RECT 1.01 0.1419 1.038 0.366 ;
        RECT 1.01 0.366 1.038 0.672 ;
        RECT 1.038 0.114 1.352 0.1419 ;
        RECT 1.352 0.114 1.3799 0.1419 ;
        RECT 1.352 0.1419 1.3799 0.366 ;
        RECT 1.106 0.638 1.3899 0.666 ;
  END
END DFFSNQ_X1

MACRO FA_X1
  CLASS core ;
  FOREIGN FA_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.536 BY 0.768 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.21 0.466 1.098 0.494 ;
      LAYER V1 ;
        RECT 0.656 0.466 0.684 0.494 ;
        RECT 1.038 0.466 1.066 0.494 ;
      LAYER M1 ;
        RECT 0.656 0.402 0.684 0.526 ;
        RECT 1.038 0.274 1.074 0.526 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.274 0.274 0.789 0.302 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.146 0.21 1.262 0.238 ;
      LAYER V1 ;
        RECT 0.178 0.21 0.206 0.238 ;
        RECT 0.58 0.21 0.608 0.238 ;
        RECT 1.202 0.21 1.23 0.238 ;
      LAYER M1 ;
        RECT 0.178 0.194 0.206 0.59 ;
        RECT 0.58 0.194 0.608 0.366 ;
        RECT 1.202 0.178 1.23 0.366 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.458 0.114 1.486 0.654 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.8179 0.207 0.846 0.64 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.1419 0.796 ;
        RECT 0.1419 0.74 0.27 0.796 ;
        RECT 0.27 0.74 0.334 0.796 ;
        RECT 0.334 0.74 0.656 0.796 ;
        RECT 0.656 0.74 0.767 0.796 ;
        RECT 0.767 0.74 1.038 0.796 ;
        RECT 1.038 0.74 1.084 0.796 ;
        RECT 1.084 0.74 1.166 0.796 ;
        RECT 1.166 0.74 1.289 0.796 ;
        RECT 1.289 0.74 1.358 0.796 ;
        RECT 1.358 0.74 1.546 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.546 0.028 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.082 0.402 1.321 0.43 ;
        RECT 0.402 0.338 1.3899 0.366 ;
      LAYER MINT1 ;
        RECT 0.082 0.402 1.321 0.43 ;
        RECT 0.402 0.338 1.3899 0.366 ;
      LAYER M1 ;
        RECT 0.027 0.178 0.065 0.338 ;
        RECT 0.027 0.338 0.065 0.366 ;
        RECT 0.065 0.338 0.103 0.366 ;
        RECT 0.103 0.338 0.1419 0.366 ;
        RECT 0.103 0.366 0.1419 0.462 ;
        RECT 0.242 0.274 0.27 0.59 ;
        RECT 0.424 0.274 0.462 0.507 ;
        RECT 0.37 0.097 0.618 0.135 ;
        RECT 0.37 0.575 0.402 0.603 ;
        RECT 0.37 0.603 0.402 0.6979 ;
        RECT 0.402 0.575 0.624 0.603 ;
        RECT 0.624 0.575 0.656 0.603 ;
        RECT 0.624 0.603 0.656 0.6979 ;
        RECT 0.624 0.6979 0.656 0.704 ;
        RECT 0.729 0.244 0.767 0.464 ;
        RECT 0.882 0.194 0.91 0.366 ;
        RECT 0.882 0.562 0.91 0.59 ;
        RECT 0.882 0.59 0.91 0.6959 ;
        RECT 0.91 0.562 1.01 0.59 ;
        RECT 1.01 0.562 1.038 0.59 ;
        RECT 1.01 0.59 1.038 0.6959 ;
        RECT 1.1379 0.072 1.166 0.6959 ;
        RECT 1.2609 0.386 1.289 0.59 ;
        RECT 0.306 0.096 0.334 0.672 ;
        RECT 0.498 0.274 0.526 0.507 ;
        RECT 0.946 0.274 0.984 0.494 ;
        RECT 0.846 0.1 1.084 0.132 ;
        RECT 1.33 0.274 1.358 0.526 ;
      LAYER V1 ;
        RECT 0.114 0.402 0.1419 0.43 ;
        RECT 0.242 0.466 0.27 0.494 ;
        RECT 0.306 0.274 0.334 0.302 ;
        RECT 0.434 0.338 0.462 0.366 ;
        RECT 0.498 0.402 0.526 0.43 ;
        RECT 0.729 0.274 0.757 0.302 ;
        RECT 0.882 0.21 0.91 0.238 ;
        RECT 0.956 0.402 0.984 0.43 ;
        RECT 1.1379 0.338 1.166 0.366 ;
        RECT 1.2609 0.402 1.289 0.43 ;
        RECT 1.33 0.338 1.358 0.366 ;
      LAYER M1 ;
        RECT 0.027 0.178 0.065 0.338 ;
        RECT 0.027 0.338 0.065 0.366 ;
        RECT 0.065 0.338 0.103 0.366 ;
        RECT 0.103 0.338 0.1419 0.366 ;
        RECT 0.103 0.366 0.1419 0.462 ;
        RECT 0.242 0.274 0.27 0.59 ;
        RECT 0.424 0.274 0.462 0.507 ;
        RECT 0.37 0.097 0.618 0.135 ;
        RECT 0.37 0.575 0.402 0.603 ;
        RECT 0.37 0.603 0.402 0.6979 ;
        RECT 0.402 0.575 0.624 0.603 ;
        RECT 0.624 0.575 0.656 0.603 ;
        RECT 0.624 0.603 0.656 0.6979 ;
        RECT 0.624 0.6979 0.656 0.704 ;
        RECT 0.729 0.244 0.767 0.464 ;
        RECT 0.882 0.194 0.91 0.366 ;
        RECT 0.882 0.562 0.91 0.59 ;
        RECT 0.882 0.59 0.91 0.6959 ;
        RECT 0.91 0.562 1.01 0.59 ;
        RECT 1.01 0.562 1.038 0.59 ;
        RECT 1.01 0.59 1.038 0.6959 ;
        RECT 1.1379 0.072 1.166 0.6959 ;
        RECT 1.2609 0.386 1.289 0.59 ;
        RECT 0.306 0.096 0.334 0.672 ;
        RECT 0.498 0.274 0.526 0.507 ;
        RECT 0.946 0.274 0.984 0.494 ;
        RECT 0.846 0.1 1.084 0.132 ;
        RECT 1.33 0.274 1.358 0.526 ;
  END
END FA_X1

MACRO FILLTIE
  CLASS core ;
  FOREIGN FILLTIE 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.578 BY 0.768 ;
  OBS
      LAYER M1 ;
        RECT -0.01 -0.028 0.588 0.028 ;
        RECT -0.01 0.74 0.588 0.796 ;
      LAYER M1 ;
        RECT -0.01 -0.028 0.588 0.028 ;
        RECT -0.01 0.74 0.588 0.796 ;
  END
END FILLTIE

MACRO FILL_X1
  CLASS core ;
  FOREIGN FILL_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.128 BY 0.768 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.138 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.138 0.028 ;
    END
  END VSS
END FILL_X1

MACRO FILL_X2
  CLASS core ;
  FOREIGN FILL_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.192 BY 0.768 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.202 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.202 0.028 ;
    END
  END VSS
END FILL_X2

MACRO FILL_X4
  CLASS core ;
  FOREIGN FILL_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.32 BY 0.768 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.33 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.33 0.028 ;
    END
  END VSS
END FILL_X4

MACRO FILL_X8
  CLASS core ;
  FOREIGN FILL_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.768 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
END FILL_X8

MACRO FILL_X16
  CLASS core ;
  FOREIGN FILL_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.088 BY 0.768 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.098 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.098 0.028 ;
    END
  END VSS
END FILL_X16

MACRO HA_X1
  CLASS core ;
  FOREIGN HA_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.832 BY 0.768 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.274 0.27 0.556 ;
        RECT 0.242 0.556 0.27 0.584 ;
        RECT 0.27 0.556 0.434 0.584 ;
        RECT 0.434 0.274 0.462 0.556 ;
        RECT 0.434 0.556 0.462 0.584 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.256 0.334 0.512 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.082 0.078 0.638 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.754 0.18 0.782 0.638 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.596 0.796 ;
        RECT 0.596 0.74 0.66 0.796 ;
        RECT 0.66 0.74 0.842 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.842 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.338 0.1019 0.622 0.13 ;
        RECT 0.406 0.184 0.498 0.216 ;
        RECT 0.498 0.184 0.53 0.216 ;
        RECT 0.498 0.216 0.53 0.462 ;
        RECT 0.498 0.462 0.53 0.602 ;
        RECT 0.53 0.184 0.632 0.216 ;
        RECT 0.632 0.184 0.66 0.216 ;
        RECT 0.632 0.216 0.66 0.462 ;
        RECT 0.114 0.166 0.1419 0.198 ;
        RECT 0.114 0.198 0.1419 0.274 ;
        RECT 0.114 0.274 0.1419 0.638 ;
        RECT 0.114 0.638 0.1419 0.666 ;
        RECT 0.1419 0.166 0.37 0.198 ;
        RECT 0.1419 0.638 0.37 0.666 ;
        RECT 0.37 0.638 0.5659 0.666 ;
        RECT 0.5659 0.274 0.596 0.638 ;
        RECT 0.5659 0.638 0.596 0.666 ;
      LAYER M1 ;
        RECT 0.338 0.1019 0.622 0.13 ;
        RECT 0.406 0.184 0.498 0.216 ;
        RECT 0.498 0.184 0.53 0.216 ;
        RECT 0.498 0.216 0.53 0.462 ;
        RECT 0.498 0.462 0.53 0.602 ;
        RECT 0.53 0.184 0.632 0.216 ;
        RECT 0.632 0.184 0.66 0.216 ;
        RECT 0.632 0.216 0.66 0.462 ;
        RECT 0.114 0.166 0.1419 0.198 ;
        RECT 0.114 0.198 0.1419 0.274 ;
        RECT 0.114 0.274 0.1419 0.638 ;
        RECT 0.114 0.638 0.1419 0.666 ;
        RECT 0.1419 0.166 0.37 0.198 ;
        RECT 0.1419 0.638 0.37 0.666 ;
        RECT 0.37 0.638 0.5659 0.666 ;
        RECT 0.5659 0.274 0.596 0.638 ;
        RECT 0.5659 0.638 0.596 0.666 ;
  END
END HA_X1

MACRO INV_X1
  CLASS core ;
  FOREIGN INV_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.192 BY 0.768 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.576 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.114 0.1419 0.64 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.202 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.202 0.028 ;
    END
  END VSS
END INV_X1

MACRO INV_X2
  CLASS core ;
  FOREIGN INV_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.256 BY 0.768 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.576 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.13 0.1419 0.576 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.266 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.266 0.028 ;
    END
  END VSS
END INV_X2

MACRO INV_X4
  CLASS core ;
  FOREIGN INV_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.768 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.048 0.256 0.08 0.368 ;
        RECT 0.048 0.368 0.08 0.396 ;
        RECT 0.048 0.396 0.08 0.512 ;
        RECT 0.08 0.368 0.238 0.396 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.041 0.1419 0.059 0.2 ;
        RECT 0.059 0.1419 0.306 0.2 ;
        RECT 0.059 0.5679 0.306 0.626 ;
        RECT 0.306 0.1419 0.334 0.2 ;
        RECT 0.306 0.2 0.334 0.5679 ;
        RECT 0.306 0.5679 0.334 0.626 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
END INV_X4

MACRO INV_X8
  CLASS core ;
  FOREIGN INV_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.64 BY 0.768 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.194 0.1419 0.396 ;
        RECT 0.114 0.396 0.1419 0.455 ;
        RECT 0.114 0.455 0.1419 0.576 ;
        RECT 0.1419 0.396 0.462 0.455 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.041 0.631 0.054 0.659 ;
        RECT 0.054 0.11 0.557 0.138 ;
        RECT 0.054 0.631 0.557 0.659 ;
        RECT 0.557 0.11 0.595 0.138 ;
        RECT 0.557 0.138 0.595 0.631 ;
        RECT 0.557 0.631 0.595 0.659 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.65 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.65 0.028 ;
    END
  END VSS
END INV_X8

MACRO INV_X12
  CLASS core ;
  FOREIGN INV_X12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.896 BY 0.768 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.192 0.1419 0.368 ;
        RECT 0.114 0.368 0.1419 0.396 ;
        RECT 0.114 0.396 0.1419 0.576 ;
        RECT 0.1419 0.368 0.686 0.396 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.054 0.1019 0.8129 0.13 ;
        RECT 0.054 0.636 0.8129 0.668 ;
        RECT 0.8129 0.1019 0.851 0.13 ;
        RECT 0.8129 0.13 0.851 0.636 ;
        RECT 0.8129 0.636 0.851 0.668 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.906 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.906 0.028 ;
    END
  END VSS
END INV_X12

MACRO INV_X16
  CLASS core ;
  FOREIGN INV_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.152 BY 0.768 ;
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.37 ;
        RECT 0.05 0.37 0.078 0.398 ;
        RECT 0.05 0.398 0.078 0.5629 ;
        RECT 0.078 0.37 0.942 0.398 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.07 0.796 ;
        RECT 1.07 0.74 1.162 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.162 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.054 0.1 1.038 0.132 ;
        RECT 0.054 0.622 1.038 0.681 ;
        RECT 1.038 0.1 1.07 0.132 ;
        RECT 1.038 0.132 1.07 0.622 ;
        RECT 1.038 0.622 1.07 0.681 ;
      LAYER M1 ;
        RECT 0.054 0.1 1.038 0.132 ;
        RECT 0.054 0.622 1.038 0.681 ;
        RECT 1.038 0.1 1.07 0.132 ;
        RECT 1.038 0.132 1.07 0.622 ;
        RECT 1.038 0.622 1.07 0.681 ;
  END
END INV_X16

MACRO LHQ_X1
  CLASS core ;
  FOREIGN LHQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.896 BY 0.768 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.16 0.27 0.512 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.512 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.8179 0.13 0.846 0.638 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.782 0.796 ;
        RECT 0.782 0.74 0.906 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.906 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.556 0.05 0.584 ;
        RECT 0.048 0.584 0.05 0.704 ;
        RECT 0.05 0.064 0.078 0.092 ;
        RECT 0.05 0.092 0.078 0.184 ;
        RECT 0.05 0.184 0.078 0.212 ;
        RECT 0.05 0.556 0.078 0.584 ;
        RECT 0.05 0.584 0.078 0.704 ;
        RECT 0.078 0.064 0.08 0.092 ;
        RECT 0.078 0.184 0.08 0.212 ;
        RECT 0.078 0.556 0.08 0.584 ;
        RECT 0.078 0.584 0.08 0.704 ;
        RECT 0.08 0.064 0.114 0.092 ;
        RECT 0.08 0.184 0.114 0.212 ;
        RECT 0.08 0.556 0.114 0.584 ;
        RECT 0.114 0.064 0.1419 0.092 ;
        RECT 0.114 0.184 0.1419 0.212 ;
        RECT 0.114 0.212 0.1419 0.322 ;
        RECT 0.114 0.322 0.1419 0.35 ;
        RECT 0.114 0.35 0.1419 0.414 ;
        RECT 0.114 0.414 0.1419 0.556 ;
        RECT 0.114 0.556 0.1419 0.584 ;
        RECT 0.1419 0.064 0.324 0.092 ;
        RECT 0.324 0.064 0.352 0.092 ;
        RECT 0.324 0.092 0.352 0.184 ;
        RECT 0.324 0.184 0.352 0.212 ;
        RECT 0.324 0.212 0.352 0.322 ;
        RECT 0.324 0.322 0.352 0.35 ;
        RECT 0.352 0.322 0.37 0.35 ;
        RECT 0.37 0.322 0.398 0.35 ;
        RECT 0.37 0.35 0.398 0.414 ;
        RECT 0.53 0.114 0.558 0.1419 ;
        RECT 0.53 0.1419 0.558 0.494 ;
        RECT 0.558 0.114 0.6899 0.1419 ;
        RECT 0.6899 0.114 0.718 0.1419 ;
        RECT 0.6899 0.1419 0.718 0.494 ;
        RECT 0.6899 0.494 0.718 0.593 ;
        RECT 0.178 0.136 0.206 0.46 ;
        RECT 0.178 0.46 0.206 0.556 ;
        RECT 0.178 0.556 0.206 0.584 ;
        RECT 0.206 0.556 0.306 0.584 ;
        RECT 0.306 0.46 0.34 0.556 ;
        RECT 0.306 0.556 0.34 0.584 ;
        RECT 0.274 0.638 0.388 0.666 ;
        RECT 0.388 0.114 0.466 0.1729 ;
        RECT 0.388 0.638 0.466 0.666 ;
        RECT 0.466 0.114 0.494 0.1729 ;
        RECT 0.466 0.1729 0.494 0.306 ;
        RECT 0.466 0.306 0.494 0.637 ;
        RECT 0.466 0.637 0.494 0.638 ;
        RECT 0.466 0.638 0.494 0.666 ;
        RECT 0.494 0.637 0.754 0.638 ;
        RECT 0.494 0.638 0.754 0.666 ;
        RECT 0.754 0.306 0.782 0.637 ;
        RECT 0.754 0.637 0.782 0.638 ;
        RECT 0.754 0.638 0.782 0.666 ;
      LAYER M1 ;
        RECT 0.048 0.556 0.05 0.584 ;
        RECT 0.048 0.584 0.05 0.704 ;
        RECT 0.05 0.064 0.078 0.092 ;
        RECT 0.05 0.092 0.078 0.184 ;
        RECT 0.05 0.184 0.078 0.212 ;
        RECT 0.05 0.556 0.078 0.584 ;
        RECT 0.05 0.584 0.078 0.704 ;
        RECT 0.078 0.064 0.08 0.092 ;
        RECT 0.078 0.184 0.08 0.212 ;
        RECT 0.078 0.556 0.08 0.584 ;
        RECT 0.078 0.584 0.08 0.704 ;
        RECT 0.08 0.064 0.114 0.092 ;
        RECT 0.08 0.184 0.114 0.212 ;
        RECT 0.08 0.556 0.114 0.584 ;
        RECT 0.114 0.064 0.1419 0.092 ;
        RECT 0.114 0.184 0.1419 0.212 ;
        RECT 0.114 0.212 0.1419 0.322 ;
        RECT 0.114 0.322 0.1419 0.35 ;
        RECT 0.114 0.35 0.1419 0.414 ;
        RECT 0.114 0.414 0.1419 0.556 ;
        RECT 0.114 0.556 0.1419 0.584 ;
        RECT 0.1419 0.064 0.324 0.092 ;
        RECT 0.324 0.064 0.352 0.092 ;
        RECT 0.324 0.092 0.352 0.184 ;
        RECT 0.324 0.184 0.352 0.212 ;
        RECT 0.324 0.212 0.352 0.322 ;
        RECT 0.324 0.322 0.352 0.35 ;
        RECT 0.352 0.322 0.37 0.35 ;
        RECT 0.37 0.322 0.398 0.35 ;
        RECT 0.37 0.35 0.398 0.414 ;
        RECT 0.53 0.114 0.558 0.1419 ;
        RECT 0.53 0.1419 0.558 0.494 ;
        RECT 0.558 0.114 0.6899 0.1419 ;
        RECT 0.6899 0.114 0.718 0.1419 ;
        RECT 0.6899 0.1419 0.718 0.494 ;
        RECT 0.6899 0.494 0.718 0.593 ;
        RECT 0.178 0.136 0.206 0.46 ;
        RECT 0.178 0.46 0.206 0.556 ;
        RECT 0.178 0.556 0.206 0.584 ;
        RECT 0.206 0.556 0.306 0.584 ;
        RECT 0.306 0.46 0.34 0.556 ;
        RECT 0.306 0.556 0.34 0.584 ;
        RECT 0.274 0.638 0.388 0.666 ;
        RECT 0.388 0.114 0.466 0.1729 ;
        RECT 0.388 0.638 0.466 0.666 ;
        RECT 0.466 0.114 0.494 0.1729 ;
        RECT 0.466 0.1729 0.494 0.306 ;
        RECT 0.466 0.306 0.494 0.637 ;
        RECT 0.466 0.637 0.494 0.638 ;
        RECT 0.466 0.638 0.494 0.666 ;
        RECT 0.494 0.637 0.754 0.638 ;
        RECT 0.494 0.638 0.754 0.666 ;
        RECT 0.754 0.306 0.782 0.637 ;
        RECT 0.754 0.637 0.782 0.638 ;
        RECT 0.754 0.638 0.782 0.666 ;
  END
END LHQ_X1

MACRO MUX2_X1
  CLASS core ;
  FOREIGN MUX2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.832 BY 0.768 ;
  PIN I0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.562 0.242 0.59 0.526 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.1419 0.448 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.118 0.658 0.394 0.686 ;
      LAYER V1 ;
        RECT 0.15 0.658 0.206 0.686 ;
      LAYER M1 ;
        RECT 0.027 0.242 0.055 0.658 ;
        RECT 0.027 0.658 0.055 0.686 ;
        RECT 0.055 0.658 0.222 0.686 ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.6899 0.192 0.718 0.638 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.462 0.796 ;
        RECT 0.462 0.74 0.526 0.796 ;
        RECT 0.526 0.74 0.782 0.796 ;
        RECT 0.782 0.74 0.842 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.842 0.028 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.274 0.338 0.558 0.366 ;
      LAYER MINT1 ;
        RECT 0.274 0.338 0.558 0.366 ;
      LAYER M1 ;
        RECT 0.08 0.162 0.099 0.19 ;
        RECT 0.099 0.162 0.157 0.19 ;
        RECT 0.099 0.492 0.157 0.52 ;
        RECT 0.099 0.52 0.157 0.576 ;
        RECT 0.157 0.162 0.306 0.19 ;
        RECT 0.157 0.492 0.306 0.52 ;
        RECT 0.306 0.162 0.334 0.19 ;
        RECT 0.306 0.19 0.334 0.492 ;
        RECT 0.306 0.492 0.334 0.52 ;
        RECT 0.29 0.658 0.434 0.704 ;
        RECT 0.434 0.306 0.462 0.658 ;
        RECT 0.434 0.658 0.462 0.704 ;
        RECT 0.498 0.274 0.526 0.428 ;
        RECT 0.37 0.0869 0.398 0.146 ;
        RECT 0.37 0.146 0.398 0.494 ;
        RECT 0.37 0.494 0.398 0.614 ;
        RECT 0.398 0.0869 0.754 0.146 ;
        RECT 0.754 0.0869 0.782 0.146 ;
        RECT 0.754 0.146 0.782 0.494 ;
      LAYER V1 ;
        RECT 0.306 0.338 0.334 0.366 ;
        RECT 0.306 0.658 0.362 0.686 ;
        RECT 0.498 0.338 0.526 0.366 ;
      LAYER M1 ;
        RECT 0.08 0.162 0.099 0.19 ;
        RECT 0.099 0.162 0.157 0.19 ;
        RECT 0.099 0.492 0.157 0.52 ;
        RECT 0.099 0.52 0.157 0.576 ;
        RECT 0.157 0.162 0.306 0.19 ;
        RECT 0.157 0.492 0.306 0.52 ;
        RECT 0.306 0.162 0.334 0.19 ;
        RECT 0.306 0.19 0.334 0.492 ;
        RECT 0.306 0.492 0.334 0.52 ;
        RECT 0.29 0.658 0.434 0.704 ;
        RECT 0.434 0.306 0.462 0.658 ;
        RECT 0.434 0.658 0.462 0.704 ;
        RECT 0.498 0.274 0.526 0.428 ;
        RECT 0.37 0.0869 0.398 0.146 ;
        RECT 0.37 0.146 0.398 0.494 ;
        RECT 0.37 0.494 0.398 0.614 ;
        RECT 0.398 0.0869 0.754 0.146 ;
        RECT 0.754 0.0869 0.782 0.146 ;
        RECT 0.754 0.146 0.782 0.494 ;
  END
END MUX2_X1

MACRO NAND2_X1
  CLASS core ;
  FOREIGN NAND2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.256 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.256 0.206 0.574 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.574 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.133 0.1419 0.192 ;
        RECT 0.114 0.192 0.1419 0.638 ;
        RECT 0.1419 0.133 0.176 0.192 ;
        RECT 0.176 0.064 0.208 0.133 ;
        RECT 0.176 0.133 0.208 0.192 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.266 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.266 0.028 ;
    END
  END VSS
END NAND2_X1

MACRO NAND2_X2
  CLASS core ;
  FOREIGN NAND2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.225 0.206 0.553 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.274 0.078 0.676 ;
        RECT 0.05 0.676 0.078 0.704 ;
        RECT 0.078 0.676 0.306 0.704 ;
        RECT 0.306 0.274 0.334 0.676 ;
        RECT 0.306 0.676 0.334 0.704 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.123 0.1419 0.181 ;
        RECT 0.114 0.181 0.1419 0.424 ;
        RECT 0.114 0.424 0.1419 0.597 ;
        RECT 0.114 0.597 0.1419 0.64 ;
        RECT 0.1419 0.123 0.242 0.181 ;
        RECT 0.1419 0.597 0.242 0.64 ;
        RECT 0.242 0.123 0.27 0.181 ;
        RECT 0.242 0.424 0.27 0.597 ;
        RECT 0.242 0.597 0.27 0.64 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
END NAND2_X2

MACRO NAND3_X1
  CLASS core ;
  FOREIGN NAND3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.32 0.27 0.448 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.255 0.206 0.512 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.215 0.078 0.574 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.082 0.1419 0.11 ;
        RECT 0.114 0.11 0.1419 0.256 ;
        RECT 0.114 0.256 0.1419 0.512 ;
        RECT 0.114 0.512 0.1419 0.676 ;
        RECT 0.114 0.676 0.1419 0.704 ;
        RECT 0.1419 0.082 0.242 0.11 ;
        RECT 0.1419 0.676 0.242 0.704 ;
        RECT 0.242 0.064 0.304 0.082 ;
        RECT 0.242 0.082 0.304 0.11 ;
        RECT 0.242 0.676 0.304 0.704 ;
        RECT 0.304 0.064 0.306 0.082 ;
        RECT 0.304 0.082 0.306 0.11 ;
        RECT 0.304 0.11 0.306 0.256 ;
        RECT 0.304 0.676 0.306 0.704 ;
        RECT 0.306 0.064 0.334 0.082 ;
        RECT 0.306 0.082 0.334 0.11 ;
        RECT 0.306 0.11 0.334 0.256 ;
        RECT 0.306 0.512 0.334 0.676 ;
        RECT 0.306 0.676 0.334 0.704 ;
        RECT 0.334 0.064 0.336 0.082 ;
        RECT 0.334 0.082 0.336 0.11 ;
        RECT 0.334 0.11 0.336 0.256 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
END NAND3_X1

MACRO NAND3_X2
  CLASS core ;
  FOREIGN NAND3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.32 0.526 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.301 0.249 0.339 0.512 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.1419 0.512 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.027 0.5679 0.366 0.626 ;
        RECT 0.366 0.5679 0.434 0.626 ;
        RECT 0.434 0.186 0.462 0.5679 ;
        RECT 0.434 0.5679 0.462 0.626 ;
        RECT 0.462 0.5679 0.494 0.626 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.366 0.796 ;
        RECT 0.366 0.74 0.526 0.796 ;
        RECT 0.526 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.21 0.111 0.498 0.1409 ;
        RECT 0.498 0.111 0.526 0.1409 ;
        RECT 0.498 0.1409 0.526 0.225 ;
        RECT 0.05 0.177 0.366 0.209 ;
      LAYER M1 ;
        RECT 0.21 0.111 0.498 0.1409 ;
        RECT 0.498 0.111 0.526 0.1409 ;
        RECT 0.498 0.1409 0.526 0.225 ;
        RECT 0.05 0.177 0.366 0.209 ;
  END
END NAND3_X2

MACRO NAND4_X1
  CLASS core ;
  FOREIGN NAND4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.448 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.256 0.398 0.574 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.242 0.27 0.512 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.194 0.206 0.448 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.194 0.078 0.574 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.512 0.1419 0.645 ;
        RECT 0.114 0.645 0.1419 0.704 ;
        RECT 0.1419 0.645 0.306 0.704 ;
        RECT 0.306 0.164 0.334 0.192 ;
        RECT 0.306 0.192 0.334 0.512 ;
        RECT 0.306 0.512 0.334 0.645 ;
        RECT 0.306 0.645 0.334 0.704 ;
        RECT 0.334 0.164 0.365 0.192 ;
        RECT 0.365 0.064 0.403 0.164 ;
        RECT 0.365 0.164 0.403 0.192 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.458 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.458 0.028 ;
    END
  END VSS
END NAND4_X1

MACRO NAND4_X2
  CLASS core ;
  FOREIGN NAND4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.704 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.358 0.594 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.34 0.398 0.526 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.242 0.206 0.512 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.257 0.078 0.512 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.112 0.555 0.144 0.576 ;
        RECT 0.112 0.576 0.144 0.638 ;
        RECT 0.112 0.638 0.144 0.666 ;
        RECT 0.144 0.638 0.434 0.666 ;
        RECT 0.434 0.294 0.462 0.322 ;
        RECT 0.434 0.322 0.462 0.548 ;
        RECT 0.434 0.548 0.462 0.555 ;
        RECT 0.434 0.555 0.462 0.576 ;
        RECT 0.434 0.638 0.462 0.666 ;
        RECT 0.462 0.294 0.562 0.322 ;
        RECT 0.462 0.548 0.562 0.555 ;
        RECT 0.462 0.555 0.562 0.576 ;
        RECT 0.462 0.638 0.562 0.666 ;
        RECT 0.562 0.294 0.59 0.322 ;
        RECT 0.562 0.548 0.59 0.555 ;
        RECT 0.562 0.555 0.59 0.576 ;
        RECT 0.562 0.576 0.59 0.638 ;
        RECT 0.562 0.638 0.59 0.666 ;
        RECT 0.59 0.294 0.654 0.322 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.656 0.796 ;
        RECT 0.656 0.74 0.714 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.714 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.1019 0.08 0.13 ;
        RECT 0.048 0.13 0.08 0.213 ;
        RECT 0.08 0.1019 0.43 0.13 ;
        RECT 0.274 0.23 0.624 0.258 ;
        RECT 0.624 0.064 0.656 0.23 ;
        RECT 0.624 0.23 0.656 0.258 ;
        RECT 0.146 0.166 0.494 0.194 ;
      LAYER M1 ;
        RECT 0.048 0.1019 0.08 0.13 ;
        RECT 0.048 0.13 0.08 0.213 ;
        RECT 0.08 0.1019 0.43 0.13 ;
        RECT 0.274 0.23 0.624 0.258 ;
        RECT 0.624 0.064 0.656 0.23 ;
        RECT 0.624 0.23 0.656 0.258 ;
        RECT 0.146 0.166 0.494 0.194 ;
  END
END NAND4_X2

MACRO NOR2_X1
  CLASS core ;
  FOREIGN NOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.256 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.194 0.206 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.194 0.078 0.512 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.13 0.1419 0.576 ;
        RECT 0.114 0.576 0.1419 0.635 ;
        RECT 0.1419 0.576 0.176 0.635 ;
        RECT 0.176 0.576 0.208 0.635 ;
        RECT 0.176 0.635 0.208 0.704 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.266 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.266 0.028 ;
    END
  END VSS
END NOR2_X1

MACRO NOR2_X2
  CLASS core ;
  FOREIGN NOR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.215 0.206 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.064 0.078 0.092 ;
        RECT 0.05 0.092 0.078 0.494 ;
        RECT 0.078 0.064 0.306 0.092 ;
        RECT 0.306 0.064 0.334 0.092 ;
        RECT 0.306 0.092 0.334 0.494 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.128 0.1419 0.156 ;
        RECT 0.114 0.156 0.1419 0.3439 ;
        RECT 0.114 0.3439 0.1419 0.556 ;
        RECT 0.114 0.556 0.1419 0.584 ;
        RECT 0.1419 0.128 0.176 0.156 ;
        RECT 0.1419 0.556 0.176 0.584 ;
        RECT 0.176 0.128 0.208 0.156 ;
        RECT 0.176 0.556 0.208 0.584 ;
        RECT 0.176 0.584 0.208 0.64 ;
        RECT 0.208 0.128 0.242 0.156 ;
        RECT 0.242 0.128 0.27 0.156 ;
        RECT 0.242 0.156 0.27 0.3439 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
END NOR2_X2

MACRO NOR3_X1
  CLASS core ;
  FOREIGN NOR3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.32 0.27 0.448 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.194 0.206 0.553 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.194 0.078 0.553 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.064 0.1419 0.092 ;
        RECT 0.114 0.092 0.1419 0.256 ;
        RECT 0.114 0.256 0.1419 0.512 ;
        RECT 0.114 0.512 0.1419 0.614 ;
        RECT 0.114 0.614 0.1419 0.642 ;
        RECT 0.1419 0.064 0.303 0.092 ;
        RECT 0.1419 0.614 0.303 0.642 ;
        RECT 0.303 0.064 0.304 0.092 ;
        RECT 0.303 0.092 0.304 0.256 ;
        RECT 0.303 0.614 0.304 0.642 ;
        RECT 0.304 0.064 0.336 0.092 ;
        RECT 0.304 0.092 0.336 0.256 ;
        RECT 0.304 0.512 0.336 0.614 ;
        RECT 0.304 0.614 0.336 0.642 ;
        RECT 0.304 0.642 0.336 0.704 ;
        RECT 0.336 0.064 0.337 0.092 ;
        RECT 0.336 0.092 0.337 0.256 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
END NOR3_X1

MACRO NOR3_X2
  CLASS core ;
  FOREIGN NOR3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.256 0.526 0.448 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.256 0.334 0.513 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.519 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.0859 0.154 0.434 0.212 ;
        RECT 0.434 0.154 0.462 0.212 ;
        RECT 0.434 0.212 0.462 0.576 ;
        RECT 0.462 0.154 0.49 0.212 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.526 0.796 ;
        RECT 0.526 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.21 0.627 0.498 0.655 ;
        RECT 0.498 0.516 0.526 0.627 ;
        RECT 0.498 0.627 0.526 0.655 ;
        RECT 0.0859 0.557 0.38 0.591 ;
      LAYER M1 ;
        RECT 0.21 0.627 0.498 0.655 ;
        RECT 0.498 0.516 0.526 0.627 ;
        RECT 0.498 0.627 0.526 0.655 ;
        RECT 0.0859 0.557 0.38 0.591 ;
  END
END NOR3_X2

MACRO NOR4_X1
  CLASS core ;
  FOREIGN NOR4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.448 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.194 0.398 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.194 0.27 0.512 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.256 0.206 0.574 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.194 0.078 0.574 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.064 0.1419 0.1019 ;
        RECT 0.114 0.1019 0.1419 0.215 ;
        RECT 0.1419 0.064 0.306 0.1019 ;
        RECT 0.306 0.064 0.334 0.1019 ;
        RECT 0.306 0.1019 0.334 0.215 ;
        RECT 0.306 0.215 0.334 0.576 ;
        RECT 0.306 0.576 0.334 0.604 ;
        RECT 0.334 0.576 0.365 0.604 ;
        RECT 0.365 0.576 0.403 0.604 ;
        RECT 0.365 0.604 0.403 0.704 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.458 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.458 0.028 ;
    END
  END VSS
END NOR4_X1

MACRO NOR4_X2
  CLASS core ;
  FOREIGN NOR4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.704 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.256 0.594 0.406 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.242 0.398 0.438 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.242 0.27 0.526 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.256 0.206 0.516 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.112 0.1019 0.144 0.13 ;
        RECT 0.112 0.13 0.144 0.192 ;
        RECT 0.112 0.192 0.144 0.213 ;
        RECT 0.144 0.1019 0.434 0.13 ;
        RECT 0.434 0.1019 0.462 0.13 ;
        RECT 0.434 0.192 0.462 0.213 ;
        RECT 0.434 0.213 0.462 0.22 ;
        RECT 0.434 0.22 0.462 0.442 ;
        RECT 0.434 0.442 0.462 0.47 ;
        RECT 0.462 0.1019 0.562 0.13 ;
        RECT 0.462 0.192 0.562 0.213 ;
        RECT 0.462 0.213 0.562 0.22 ;
        RECT 0.462 0.442 0.562 0.47 ;
        RECT 0.562 0.1019 0.59 0.13 ;
        RECT 0.562 0.13 0.59 0.192 ;
        RECT 0.562 0.192 0.59 0.213 ;
        RECT 0.562 0.213 0.59 0.22 ;
        RECT 0.562 0.442 0.59 0.47 ;
        RECT 0.59 0.442 0.663 0.47 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.43 0.796 ;
        RECT 0.43 0.74 0.494 0.796 ;
        RECT 0.494 0.74 0.656 0.796 ;
        RECT 0.656 0.74 0.714 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.714 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.21 0.5699 0.494 0.602 ;
        RECT 0.048 0.555 0.08 0.638 ;
        RECT 0.048 0.638 0.08 0.666 ;
        RECT 0.08 0.638 0.43 0.666 ;
        RECT 0.338 0.506 0.624 0.534 ;
        RECT 0.624 0.506 0.656 0.534 ;
        RECT 0.624 0.534 0.656 0.686 ;
      LAYER M1 ;
        RECT 0.21 0.5699 0.494 0.602 ;
        RECT 0.048 0.555 0.08 0.638 ;
        RECT 0.048 0.638 0.08 0.666 ;
        RECT 0.08 0.638 0.43 0.666 ;
        RECT 0.338 0.506 0.624 0.534 ;
        RECT 0.624 0.506 0.656 0.534 ;
        RECT 0.624 0.534 0.656 0.686 ;
  END
END NOR4_X2

MACRO OAI21_X1
  CLASS core ;
  FOREIGN OAI21_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.256 0.206 0.576 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.634 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.256 0.334 0.576 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.1419 0.636 ;
        RECT 0.114 0.636 0.1419 0.668 ;
        RECT 0.1419 0.636 0.298 0.668 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.298 0.796 ;
        RECT 0.298 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.073 0.078 0.155 ;
        RECT 0.05 0.155 0.078 0.187 ;
        RECT 0.078 0.155 0.298 0.187 ;
      LAYER M1 ;
        RECT 0.05 0.073 0.078 0.155 ;
        RECT 0.05 0.155 0.078 0.187 ;
        RECT 0.078 0.155 0.298 0.187 ;
  END
END OAI21_X1

MACRO OAI21_X2
  CLASS core ;
  FOREIGN OAI21_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.365 0.32 0.403 0.448 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.242 0.27 0.2829 ;
        RECT 0.242 0.2829 0.27 0.502 ;
        RECT 0.242 0.502 0.27 0.53 ;
        RECT 0.27 0.502 0.498 0.53 ;
        RECT 0.498 0.2829 0.526 0.502 ;
        RECT 0.498 0.502 0.526 0.53 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.256 0.1419 0.525 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.029 0.5699 0.178 0.602 ;
        RECT 0.178 0.166 0.206 0.194 ;
        RECT 0.178 0.194 0.206 0.278 ;
        RECT 0.178 0.278 0.206 0.5699 ;
        RECT 0.178 0.5699 0.206 0.602 ;
        RECT 0.206 0.166 0.426 0.194 ;
        RECT 0.206 0.5699 0.426 0.602 ;
        RECT 0.426 0.166 0.434 0.194 ;
        RECT 0.434 0.166 0.462 0.194 ;
        RECT 0.434 0.194 0.462 0.278 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.535 0.796 ;
        RECT 0.535 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.048 0.1019 0.08 0.13 ;
        RECT 0.048 0.13 0.08 0.213 ;
        RECT 0.08 0.1019 0.498 0.13 ;
        RECT 0.498 0.1019 0.526 0.13 ;
        RECT 0.498 0.13 0.526 0.213 ;
        RECT 0.498 0.213 0.526 0.215 ;
        RECT 0.146 0.638 0.535 0.666 ;
      LAYER M1 ;
        RECT 0.048 0.1019 0.08 0.13 ;
        RECT 0.048 0.13 0.08 0.213 ;
        RECT 0.08 0.1019 0.498 0.13 ;
        RECT 0.498 0.1019 0.526 0.13 ;
        RECT 0.498 0.13 0.526 0.213 ;
        RECT 0.498 0.213 0.526 0.215 ;
        RECT 0.146 0.638 0.535 0.666 ;
  END
END OAI21_X2

MACRO OAI22_X1
  CLASS core ;
  FOREIGN OAI22_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.448 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.199 0.27 0.576 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.279 0.398 0.576 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.192 0.206 0.512 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.048 0.192 0.08 0.576 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.1409 0.638 0.306 0.666 ;
        RECT 0.306 0.182 0.334 0.638 ;
        RECT 0.306 0.638 0.334 0.666 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.398 0.796 ;
        RECT 0.398 0.74 0.458 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.458 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.101 0.37 0.131 ;
        RECT 0.37 0.101 0.398 0.131 ;
        RECT 0.37 0.131 0.398 0.211 ;
      LAYER M1 ;
        RECT 0.05 0.101 0.37 0.131 ;
        RECT 0.37 0.101 0.398 0.131 ;
        RECT 0.37 0.131 0.398 0.211 ;
  END
END OAI22_X1

MACRO OAI22_X2
  CLASS core ;
  FOREIGN OAI22_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.768 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.256 0.462 0.279 ;
        RECT 0.434 0.279 0.462 0.466 ;
        RECT 0.434 0.466 0.462 0.494 ;
        RECT 0.462 0.466 0.6899 0.494 ;
        RECT 0.6899 0.279 0.718 0.466 ;
        RECT 0.6899 0.466 0.718 0.494 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.562 0.256 0.59 0.398 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.242 0.334 0.486 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.242 0.1419 0.512 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.386 0.27 0.53 ;
        RECT 0.242 0.53 0.27 0.558 ;
        RECT 0.27 0.53 0.37 0.558 ;
        RECT 0.37 0.169 0.398 0.197 ;
        RECT 0.37 0.197 0.398 0.278 ;
        RECT 0.37 0.278 0.398 0.386 ;
        RECT 0.37 0.386 0.398 0.53 ;
        RECT 0.37 0.53 0.398 0.558 ;
        RECT 0.398 0.169 0.626 0.197 ;
        RECT 0.398 0.53 0.626 0.558 ;
        RECT 0.626 0.169 0.654 0.197 ;
        RECT 0.626 0.197 0.654 0.278 ;
        RECT 0.626 0.53 0.654 0.558 ;
        RECT 0.654 0.53 0.6899 0.558 ;
        RECT 0.6899 0.53 0.718 0.558 ;
        RECT 0.6899 0.558 0.718 0.672 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.362 0.796 ;
        RECT 0.362 0.74 0.654 0.796 ;
        RECT 0.654 0.74 0.718 0.796 ;
        RECT 0.718 0.74 0.778 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.778 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.402 0.604 0.626 0.636 ;
        RECT 0.626 0.604 0.654 0.636 ;
        RECT 0.626 0.636 0.654 0.6959 ;
        RECT 0.041 0.099 0.6899 0.133 ;
        RECT 0.6899 0.099 0.718 0.133 ;
        RECT 0.6899 0.133 0.718 0.211 ;
        RECT 0.05 0.612 0.362 0.67 ;
      LAYER M1 ;
        RECT 0.402 0.604 0.626 0.636 ;
        RECT 0.626 0.604 0.654 0.636 ;
        RECT 0.626 0.636 0.654 0.6959 ;
        RECT 0.041 0.099 0.6899 0.133 ;
        RECT 0.6899 0.099 0.718 0.133 ;
        RECT 0.6899 0.133 0.718 0.211 ;
        RECT 0.05 0.612 0.362 0.67 ;
  END
END OAI22_X2

MACRO OR2_X1
  CLASS core ;
  FOREIGN OR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.384 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.096 0.206 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.243 0.078 0.641 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.114 0.334 0.64 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.27 0.796 ;
        RECT 0.27 0.74 0.394 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.394 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.13 0.1419 0.336 ;
        RECT 0.114 0.336 0.1419 0.556 ;
        RECT 0.114 0.556 0.1419 0.584 ;
        RECT 0.1419 0.556 0.242 0.584 ;
        RECT 0.242 0.336 0.27 0.556 ;
        RECT 0.242 0.556 0.27 0.584 ;
      LAYER M1 ;
        RECT 0.114 0.13 0.1419 0.336 ;
        RECT 0.114 0.336 0.1419 0.556 ;
        RECT 0.114 0.556 0.1419 0.584 ;
        RECT 0.1419 0.556 0.242 0.584 ;
        RECT 0.242 0.336 0.27 0.556 ;
        RECT 0.242 0.556 0.27 0.584 ;
  END
END OR2_X1

MACRO OR2_X2
  CLASS core ;
  FOREIGN OR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.448 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.242 0.1419 0.512 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.512 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.302 0.064 0.306 0.135 ;
        RECT 0.302 0.638 0.306 0.704 ;
        RECT 0.306 0.064 0.334 0.135 ;
        RECT 0.306 0.135 0.334 0.638 ;
        RECT 0.306 0.638 0.334 0.704 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.27 0.796 ;
        RECT 0.27 0.74 0.458 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.458 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.077 0.154 0.146 0.188 ;
        RECT 0.146 0.154 0.242 0.188 ;
        RECT 0.146 0.58 0.242 0.608 ;
        RECT 0.242 0.154 0.27 0.188 ;
        RECT 0.242 0.188 0.27 0.58 ;
        RECT 0.242 0.58 0.27 0.608 ;
      LAYER M1 ;
        RECT 0.077 0.154 0.146 0.188 ;
        RECT 0.146 0.154 0.242 0.188 ;
        RECT 0.146 0.58 0.242 0.608 ;
        RECT 0.242 0.154 0.27 0.188 ;
        RECT 0.242 0.188 0.27 0.58 ;
        RECT 0.242 0.58 0.27 0.608 ;
  END
END OR2_X2

MACRO OR3_X1
  CLASS core ;
  FOREIGN OR3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.192 0.334 0.576 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.176 0.192 0.208 0.576 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.045 0.192 0.083 0.576 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.114 0.462 0.654 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.234 0.796 ;
        RECT 0.234 0.74 0.398 0.796 ;
        RECT 0.398 0.74 0.522 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.522 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.054 0.109 0.278 0.137 ;
        RECT 0.278 0.109 0.37 0.137 ;
        RECT 0.278 0.631 0.37 0.673 ;
        RECT 0.37 0.109 0.398 0.137 ;
        RECT 0.37 0.137 0.398 0.631 ;
        RECT 0.37 0.631 0.398 0.673 ;
        RECT 0.0859 0.636 0.234 0.668 ;
      LAYER M1 ;
        RECT 0.054 0.109 0.278 0.137 ;
        RECT 0.278 0.109 0.37 0.137 ;
        RECT 0.278 0.631 0.37 0.673 ;
        RECT 0.37 0.109 0.398 0.137 ;
        RECT 0.37 0.137 0.398 0.631 ;
        RECT 0.37 0.631 0.398 0.673 ;
        RECT 0.0859 0.636 0.234 0.668 ;
  END
END OR3_X1

MACRO OR3_X2
  CLASS core ;
  FOREIGN OR3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.512 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.255 0.1419 0.448 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.256 0.078 0.526 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.231 0.27 0.448 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.366 0.064 0.37 0.13 ;
        RECT 0.366 0.636 0.37 0.704 ;
        RECT 0.37 0.064 0.398 0.13 ;
        RECT 0.37 0.13 0.398 0.636 ;
        RECT 0.37 0.636 0.398 0.704 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.302 0.796 ;
        RECT 0.302 0.74 0.334 0.796 ;
        RECT 0.334 0.74 0.522 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.522 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.5729 0.078 0.603 ;
        RECT 0.05 0.603 0.078 0.686 ;
        RECT 0.078 0.5729 0.302 0.603 ;
        RECT 0.06 0.155 0.1409 0.187 ;
        RECT 0.1409 0.155 0.306 0.187 ;
        RECT 0.1409 0.505 0.306 0.537 ;
        RECT 0.306 0.155 0.334 0.187 ;
        RECT 0.306 0.187 0.334 0.505 ;
        RECT 0.306 0.505 0.334 0.537 ;
      LAYER M1 ;
        RECT 0.05 0.5729 0.078 0.603 ;
        RECT 0.05 0.603 0.078 0.686 ;
        RECT 0.078 0.5729 0.302 0.603 ;
        RECT 0.06 0.155 0.1409 0.187 ;
        RECT 0.1409 0.155 0.306 0.187 ;
        RECT 0.1409 0.505 0.306 0.537 ;
        RECT 0.306 0.155 0.334 0.187 ;
        RECT 0.306 0.187 0.334 0.505 ;
        RECT 0.306 0.505 0.334 0.537 ;
  END
END OR3_X2

MACRO OR4_X1
  CLASS core ;
  FOREIGN OR4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.192 0.398 0.576 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.24 0.192 0.272 0.576 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.198 0.1419 0.576 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.192 0.078 0.576 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.114 0.526 0.64 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.298 0.796 ;
        RECT 0.298 0.74 0.462 0.796 ;
        RECT 0.462 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.054 0.1019 0.338 0.13 ;
        RECT 0.338 0.1019 0.434 0.13 ;
        RECT 0.338 0.63 0.434 0.662 ;
        RECT 0.434 0.1019 0.462 0.13 ;
        RECT 0.434 0.13 0.462 0.63 ;
        RECT 0.434 0.63 0.462 0.662 ;
        RECT 0.146 0.617 0.298 0.655 ;
      LAYER M1 ;
        RECT 0.054 0.1019 0.338 0.13 ;
        RECT 0.338 0.1019 0.434 0.13 ;
        RECT 0.338 0.63 0.434 0.662 ;
        RECT 0.434 0.1019 0.462 0.13 ;
        RECT 0.434 0.13 0.462 0.63 ;
        RECT 0.434 0.63 0.462 0.662 ;
        RECT 0.146 0.617 0.298 0.655 ;
  END
END OR4_X1

MACRO OR4_X2
  CLASS core ;
  FOREIGN OR4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.64 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.192 0.334 0.53 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.213 0.27 0.576 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.213 0.1419 0.576 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.191 0.078 0.576 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.496 0.128 0.528 0.704 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.302 0.796 ;
        RECT 0.302 0.74 0.46 0.796 ;
        RECT 0.46 0.74 0.65 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.65 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.146 0.623 0.302 0.681 ;
        RECT 0.054 0.0869 0.342 0.145 ;
        RECT 0.342 0.0869 0.432 0.145 ;
        RECT 0.342 0.5679 0.432 0.624 ;
        RECT 0.432 0.0869 0.46 0.145 ;
        RECT 0.432 0.145 0.46 0.5679 ;
        RECT 0.432 0.5679 0.46 0.624 ;
      LAYER M1 ;
        RECT 0.146 0.623 0.302 0.681 ;
        RECT 0.054 0.0869 0.342 0.145 ;
        RECT 0.342 0.0869 0.432 0.145 ;
        RECT 0.342 0.5679 0.432 0.624 ;
        RECT 0.432 0.0869 0.46 0.145 ;
        RECT 0.432 0.145 0.46 0.5679 ;
        RECT 0.432 0.5679 0.46 0.624 ;
  END
END OR4_X2

MACRO SDFFRNQ_X1
  CLASS core ;
  FOREIGN SDFFRNQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.92 BY 0.768 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.363 0.515 0.528 ;
        RECT 0.515 0.363 0.526 0.528 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.965 0.338 1.454 0.366 ;
        RECT 1.454 0.338 1.592 0.366 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.372 0.334 0.5719 ;
        RECT 0.306 0.5719 0.334 0.6 ;
        RECT 0.334 0.5719 0.515 0.6 ;
        RECT 0.515 0.5719 0.562 0.6 ;
        RECT 0.562 0.314 0.59 0.372 ;
        RECT 0.562 0.372 0.59 0.5719 ;
        RECT 0.562 0.5719 0.59 0.6 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.363 0.398 0.512 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.276 0.078 0.534 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.84 0.064 1.872 0.704 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.1419 0.796 ;
        RECT 0.1419 0.74 0.206 0.796 ;
        RECT 0.206 0.74 0.754 0.796 ;
        RECT 0.754 0.74 0.782 0.796 ;
        RECT 0.782 0.74 1.066 0.796 ;
        RECT 1.066 0.74 1.422 0.796 ;
        RECT 1.422 0.74 1.49 0.796 ;
        RECT 1.49 0.74 1.742 0.796 ;
        RECT 1.742 0.74 1.93 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.93 0.028 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.146 0.53 1.326 0.558 ;
        RECT 0.722 0.402 1.121 0.43 ;
        RECT 0.082 0.274 1.454 0.302 ;
      LAYER MINT1 ;
        RECT 0.146 0.53 1.326 0.558 ;
        RECT 0.722 0.402 1.121 0.43 ;
        RECT 0.082 0.274 1.454 0.302 ;
      LAYER M1 ;
        RECT 0.045 0.096 0.083 0.2039 ;
        RECT 0.045 0.2039 0.083 0.232 ;
        RECT 0.045 0.604 0.083 0.632 ;
        RECT 0.045 0.632 0.083 0.6879 ;
        RECT 0.083 0.2039 0.114 0.232 ;
        RECT 0.083 0.604 0.114 0.632 ;
        RECT 0.114 0.2039 0.1419 0.232 ;
        RECT 0.114 0.232 0.1419 0.604 ;
        RECT 0.114 0.604 0.1419 0.632 ;
        RECT 0.242 0.096 0.27 0.267 ;
        RECT 0.242 0.267 0.27 0.295 ;
        RECT 0.242 0.295 0.27 0.672 ;
        RECT 0.27 0.267 0.515 0.295 ;
        RECT 0.338 0.184 0.626 0.212 ;
        RECT 0.626 0.184 0.654 0.212 ;
        RECT 0.626 0.212 0.654 0.276 ;
        RECT 0.392 0.636 0.754 0.668 ;
        RECT 0.754 0.247 0.782 0.546 ;
        RECT 0.466 0.1019 0.878 0.13 ;
        RECT 1.061 0.24 1.098 0.446 ;
        RECT 1.202 0.171 1.23 0.511 ;
        RECT 1.458 0.146 1.49 0.6979 ;
        RECT 1.165 0.618 1.33 0.646 ;
        RECT 1.33 0.064 1.358 0.092 ;
        RECT 1.33 0.092 1.358 0.366 ;
        RECT 1.33 0.366 1.358 0.618 ;
        RECT 1.33 0.618 1.358 0.646 ;
        RECT 1.358 0.064 1.607 0.092 ;
        RECT 1.607 0.064 1.635 0.092 ;
        RECT 1.607 0.092 1.635 0.366 ;
        RECT 1.554 0.46 1.582 0.624 ;
        RECT 1.554 0.624 1.582 0.68 ;
        RECT 1.582 0.624 1.714 0.68 ;
        RECT 1.714 0.072 1.742 0.46 ;
        RECT 1.714 0.46 1.742 0.624 ;
        RECT 1.714 0.624 1.742 0.68 ;
        RECT 0.178 0.125 0.206 0.574 ;
        RECT 0.6899 0.387 0.718 0.59 ;
        RECT 0.8179 0.257 0.85 0.469 ;
        RECT 0.6899 0.166 0.718 0.194 ;
        RECT 0.6899 0.194 0.718 0.276 ;
        RECT 0.718 0.166 0.942 0.194 ;
        RECT 0.991 0.242 1.025 0.422 ;
        RECT 0.79 0.636 1.066 0.668 ;
        RECT 0.904 0.274 0.932 0.49 ;
        RECT 0.904 0.49 0.932 0.518 ;
        RECT 0.932 0.49 1.1339 0.518 ;
        RECT 1.1339 0.082 1.166 0.274 ;
        RECT 1.1339 0.274 1.166 0.49 ;
        RECT 1.1339 0.49 1.166 0.518 ;
        RECT 1.266 0.178 1.294 0.574 ;
        RECT 1.3939 0.178 1.422 0.494 ;
        RECT 1.532 0.154 1.571 0.416 ;
      LAYER V1 ;
        RECT 0.114 0.274 0.1419 0.302 ;
        RECT 0.178 0.53 0.206 0.558 ;
        RECT 0.6899 0.53 0.718 0.558 ;
        RECT 0.754 0.402 0.782 0.43 ;
        RECT 0.8179 0.274 0.846 0.302 ;
        RECT 0.997 0.338 1.025 0.366 ;
        RECT 1.061 0.402 1.089 0.43 ;
        RECT 1.202 0.274 1.23 0.302 ;
        RECT 1.266 0.53 1.294 0.558 ;
        RECT 1.3939 0.274 1.422 0.302 ;
        RECT 1.532 0.338 1.56 0.366 ;
      LAYER M1 ;
        RECT 0.045 0.096 0.083 0.2039 ;
        RECT 0.045 0.2039 0.083 0.232 ;
        RECT 0.045 0.604 0.083 0.632 ;
        RECT 0.045 0.632 0.083 0.6879 ;
        RECT 0.083 0.2039 0.114 0.232 ;
        RECT 0.083 0.604 0.114 0.632 ;
        RECT 0.114 0.2039 0.1419 0.232 ;
        RECT 0.114 0.232 0.1419 0.604 ;
        RECT 0.114 0.604 0.1419 0.632 ;
        RECT 0.242 0.096 0.27 0.267 ;
        RECT 0.242 0.267 0.27 0.295 ;
        RECT 0.242 0.295 0.27 0.672 ;
        RECT 0.27 0.267 0.515 0.295 ;
        RECT 0.338 0.184 0.626 0.212 ;
        RECT 0.626 0.184 0.654 0.212 ;
        RECT 0.626 0.212 0.654 0.276 ;
        RECT 0.392 0.636 0.754 0.668 ;
        RECT 0.754 0.247 0.782 0.546 ;
        RECT 0.466 0.1019 0.878 0.13 ;
        RECT 1.061 0.24 1.098 0.446 ;
        RECT 1.202 0.171 1.23 0.511 ;
        RECT 1.458 0.146 1.49 0.6979 ;
        RECT 1.165 0.618 1.33 0.646 ;
        RECT 1.33 0.064 1.358 0.092 ;
        RECT 1.33 0.092 1.358 0.366 ;
        RECT 1.33 0.366 1.358 0.618 ;
        RECT 1.33 0.618 1.358 0.646 ;
        RECT 1.358 0.064 1.607 0.092 ;
        RECT 1.607 0.064 1.635 0.092 ;
        RECT 1.607 0.092 1.635 0.366 ;
        RECT 1.554 0.46 1.582 0.624 ;
        RECT 1.554 0.624 1.582 0.68 ;
        RECT 1.582 0.624 1.714 0.68 ;
        RECT 1.714 0.072 1.742 0.46 ;
        RECT 1.714 0.46 1.742 0.624 ;
        RECT 1.714 0.624 1.742 0.68 ;
        RECT 0.178 0.125 0.206 0.574 ;
        RECT 0.6899 0.387 0.718 0.59 ;
        RECT 0.8179 0.257 0.85 0.469 ;
        RECT 0.6899 0.166 0.718 0.194 ;
        RECT 0.6899 0.194 0.718 0.276 ;
        RECT 0.718 0.166 0.942 0.194 ;
        RECT 0.991 0.242 1.025 0.422 ;
        RECT 0.79 0.636 1.066 0.668 ;
        RECT 0.904 0.274 0.932 0.49 ;
        RECT 0.904 0.49 0.932 0.518 ;
        RECT 0.932 0.49 1.1339 0.518 ;
        RECT 1.1339 0.082 1.166 0.274 ;
        RECT 1.1339 0.274 1.166 0.49 ;
        RECT 1.1339 0.49 1.166 0.518 ;
        RECT 1.266 0.178 1.294 0.574 ;
        RECT 1.3939 0.178 1.422 0.494 ;
        RECT 1.532 0.154 1.571 0.416 ;
  END
END SDFFRNQ_X1

MACRO SDFFSNQ_X1
  CLASS core ;
  FOREIGN SDFFSNQ_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.92 BY 0.768 ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.384 0.51 0.528 ;
        RECT 0.51 0.384 0.526 0.528 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.306 0.372 0.334 0.5719 ;
        RECT 0.306 0.5719 0.334 0.6 ;
        RECT 0.334 0.5719 0.51 0.6 ;
        RECT 0.51 0.5719 0.562 0.6 ;
        RECT 0.562 0.314 0.59 0.372 ;
        RECT 0.562 0.372 0.59 0.5719 ;
        RECT 0.562 0.5719 0.59 0.6 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.37 0.363 0.398 0.512 ;
    END
  END SI
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER MINT1 ;
        RECT 0.958 0.338 1.454 0.366 ;
        RECT 1.454 0.338 1.586 0.366 ;
    END
  END SN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.272 0.078 0.512 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.84 0.064 1.872 0.704 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.1419 0.796 ;
        RECT 0.1419 0.74 0.206 0.796 ;
        RECT 0.206 0.74 0.746 0.796 ;
        RECT 0.746 0.74 0.782 0.796 ;
        RECT 0.782 0.74 0.862 0.796 ;
        RECT 0.862 0.74 1.646 0.796 ;
        RECT 1.646 0.74 1.742 0.796 ;
        RECT 1.742 0.74 1.93 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.93 0.028 ;
    END
  END VSS
  OBS
      LAYER MINT1 ;
        RECT 0.146 0.53 1.326 0.558 ;
        RECT 0.722 0.402 1.114 0.43 ;
        RECT 0.082 0.274 1.454 0.302 ;
      LAYER MINT1 ;
        RECT 0.146 0.53 1.326 0.558 ;
        RECT 0.722 0.402 1.114 0.43 ;
        RECT 0.082 0.274 1.454 0.302 ;
      LAYER M1 ;
        RECT 0.048 0.064 0.08 0.2 ;
        RECT 0.048 0.2 0.08 0.228 ;
        RECT 0.048 0.604 0.08 0.632 ;
        RECT 0.048 0.632 0.08 0.6879 ;
        RECT 0.08 0.2 0.114 0.228 ;
        RECT 0.08 0.604 0.114 0.632 ;
        RECT 0.114 0.2 0.1419 0.228 ;
        RECT 0.114 0.228 0.1419 0.604 ;
        RECT 0.114 0.604 0.1419 0.632 ;
        RECT 0.242 0.082 0.27 0.266 ;
        RECT 0.242 0.266 0.27 0.295 ;
        RECT 0.242 0.295 0.27 0.296 ;
        RECT 0.242 0.296 0.27 0.686 ;
        RECT 0.27 0.266 0.434 0.295 ;
        RECT 0.434 0.266 0.51 0.295 ;
        RECT 0.434 0.295 0.51 0.296 ;
        RECT 0.338 0.184 0.626 0.212 ;
        RECT 0.626 0.184 0.654 0.212 ;
        RECT 0.626 0.212 0.654 0.276 ;
        RECT 0.392 0.636 0.746 0.668 ;
        RECT 0.754 0.238 0.782 0.547 ;
        RECT 0.466 0.1019 0.878 0.13 ;
        RECT 0.98 0.322 1.018 0.419 ;
        RECT 0.898 0.274 0.926 0.487 ;
        RECT 0.898 0.487 0.926 0.515 ;
        RECT 0.926 0.487 1.008 0.515 ;
        RECT 1.008 0.487 1.04 0.515 ;
        RECT 1.008 0.515 1.04 0.704 ;
        RECT 1.04 0.487 1.1379 0.515 ;
        RECT 1.1379 0.098 1.166 0.274 ;
        RECT 1.1379 0.274 1.166 0.487 ;
        RECT 1.1379 0.487 1.166 0.515 ;
        RECT 1.266 0.178 1.294 0.574 ;
        RECT 1.3939 0.178 1.422 0.402 ;
        RECT 1.526 0.184 1.554 0.403 ;
        RECT 1.402 0.638 1.646 0.666 ;
        RECT 0.178 0.096 0.206 0.619 ;
        RECT 0.654 0.387 0.682 0.574 ;
        RECT 0.83 0.257 0.862 0.469 ;
        RECT 0.6899 0.166 0.718 0.194 ;
        RECT 0.6899 0.194 0.718 0.276 ;
        RECT 0.718 0.166 0.942 0.194 ;
        RECT 1.054 0.24 1.092 0.446 ;
        RECT 1.202 0.171 1.23 0.383 ;
        RECT 1.165 0.618 1.33 0.646 ;
        RECT 1.33 0.082 1.358 0.11 ;
        RECT 1.33 0.11 1.358 0.366 ;
        RECT 1.33 0.366 1.358 0.618 ;
        RECT 1.33 0.618 1.358 0.646 ;
        RECT 1.358 0.082 1.607 0.11 ;
        RECT 1.607 0.082 1.645 0.11 ;
        RECT 1.607 0.11 1.645 0.366 ;
        RECT 1.462 0.402 1.49 0.574 ;
        RECT 1.462 0.574 1.49 0.602 ;
        RECT 1.49 0.574 1.714 0.602 ;
        RECT 1.714 0.096 1.742 0.402 ;
        RECT 1.714 0.402 1.742 0.574 ;
        RECT 1.714 0.574 1.742 0.602 ;
      LAYER V1 ;
        RECT 0.114 0.274 0.1419 0.302 ;
        RECT 0.178 0.53 0.206 0.558 ;
        RECT 0.654 0.53 0.682 0.558 ;
        RECT 0.754 0.402 0.782 0.43 ;
        RECT 0.834 0.274 0.862 0.302 ;
        RECT 0.99 0.338 1.018 0.366 ;
        RECT 1.054 0.402 1.082 0.43 ;
        RECT 1.202 0.274 1.23 0.302 ;
        RECT 1.266 0.53 1.294 0.558 ;
        RECT 1.3939 0.274 1.422 0.302 ;
        RECT 1.526 0.338 1.554 0.366 ;
      LAYER M1 ;
        RECT 0.048 0.064 0.08 0.2 ;
        RECT 0.048 0.2 0.08 0.228 ;
        RECT 0.048 0.604 0.08 0.632 ;
        RECT 0.048 0.632 0.08 0.6879 ;
        RECT 0.08 0.2 0.114 0.228 ;
        RECT 0.08 0.604 0.114 0.632 ;
        RECT 0.114 0.2 0.1419 0.228 ;
        RECT 0.114 0.228 0.1419 0.604 ;
        RECT 0.114 0.604 0.1419 0.632 ;
        RECT 0.242 0.082 0.27 0.266 ;
        RECT 0.242 0.266 0.27 0.295 ;
        RECT 0.242 0.295 0.27 0.296 ;
        RECT 0.242 0.296 0.27 0.686 ;
        RECT 0.27 0.266 0.434 0.295 ;
        RECT 0.434 0.266 0.51 0.295 ;
        RECT 0.434 0.295 0.51 0.296 ;
        RECT 0.338 0.184 0.626 0.212 ;
        RECT 0.626 0.184 0.654 0.212 ;
        RECT 0.626 0.212 0.654 0.276 ;
        RECT 0.392 0.636 0.746 0.668 ;
        RECT 0.754 0.238 0.782 0.547 ;
        RECT 0.466 0.1019 0.878 0.13 ;
        RECT 0.98 0.322 1.018 0.419 ;
        RECT 0.898 0.274 0.926 0.487 ;
        RECT 0.898 0.487 0.926 0.515 ;
        RECT 0.926 0.487 1.008 0.515 ;
        RECT 1.008 0.487 1.04 0.515 ;
        RECT 1.008 0.515 1.04 0.704 ;
        RECT 1.04 0.487 1.1379 0.515 ;
        RECT 1.1379 0.098 1.166 0.274 ;
        RECT 1.1379 0.274 1.166 0.487 ;
        RECT 1.1379 0.487 1.166 0.515 ;
        RECT 1.266 0.178 1.294 0.574 ;
        RECT 1.3939 0.178 1.422 0.402 ;
        RECT 1.526 0.184 1.554 0.403 ;
        RECT 1.402 0.638 1.646 0.666 ;
        RECT 0.178 0.096 0.206 0.619 ;
        RECT 0.654 0.387 0.682 0.574 ;
        RECT 0.83 0.257 0.862 0.469 ;
        RECT 0.6899 0.166 0.718 0.194 ;
        RECT 0.6899 0.194 0.718 0.276 ;
        RECT 0.718 0.166 0.942 0.194 ;
        RECT 1.054 0.24 1.092 0.446 ;
        RECT 1.202 0.171 1.23 0.383 ;
        RECT 1.165 0.618 1.33 0.646 ;
        RECT 1.33 0.082 1.358 0.11 ;
        RECT 1.33 0.11 1.358 0.366 ;
        RECT 1.33 0.366 1.358 0.618 ;
        RECT 1.33 0.618 1.358 0.646 ;
        RECT 1.358 0.082 1.607 0.11 ;
        RECT 1.607 0.082 1.645 0.11 ;
        RECT 1.607 0.11 1.645 0.366 ;
        RECT 1.462 0.402 1.49 0.574 ;
        RECT 1.462 0.574 1.49 0.602 ;
        RECT 1.49 0.574 1.714 0.602 ;
        RECT 1.714 0.096 1.742 0.402 ;
        RECT 1.714 0.402 1.742 0.574 ;
        RECT 1.714 0.574 1.742 0.602 ;
  END
END SDFFSNQ_X1

MACRO TBUF_X1
  CLASS core ;
  FOREIGN TBUF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.704 BY 0.768 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.384 0.1419 0.492 ;
        RECT 0.114 0.492 0.1419 0.52 ;
        RECT 0.1419 0.492 0.206 0.52 ;
        RECT 0.206 0.492 0.242 0.52 ;
        RECT 0.242 0.306 0.27 0.384 ;
        RECT 0.242 0.384 0.27 0.492 ;
        RECT 0.242 0.492 0.27 0.52 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.37 0.462 0.576 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.624 0.064 0.656 0.704 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.588 0.796 ;
        RECT 0.588 0.74 0.714 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.714 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.072 0.078 0.312 ;
        RECT 0.05 0.312 0.078 0.34 ;
        RECT 0.05 0.34 0.078 0.418 ;
        RECT 0.05 0.418 0.078 0.686 ;
        RECT 0.078 0.312 0.178 0.34 ;
        RECT 0.178 0.312 0.206 0.34 ;
        RECT 0.178 0.34 0.206 0.418 ;
        RECT 0.146 0.574 0.202 0.602 ;
        RECT 0.202 0.1019 0.23 0.13 ;
        RECT 0.202 0.13 0.23 0.23 ;
        RECT 0.202 0.23 0.23 0.258 ;
        RECT 0.202 0.574 0.23 0.602 ;
        RECT 0.23 0.1019 0.306 0.13 ;
        RECT 0.23 0.23 0.306 0.258 ;
        RECT 0.23 0.574 0.306 0.602 ;
        RECT 0.306 0.1019 0.334 0.13 ;
        RECT 0.306 0.23 0.334 0.258 ;
        RECT 0.306 0.258 0.334 0.314 ;
        RECT 0.306 0.314 0.334 0.574 ;
        RECT 0.306 0.574 0.334 0.602 ;
        RECT 0.334 0.1019 0.51 0.13 ;
        RECT 0.51 0.1019 0.542 0.13 ;
        RECT 0.51 0.13 0.542 0.23 ;
        RECT 0.51 0.23 0.542 0.258 ;
        RECT 0.51 0.258 0.542 0.314 ;
        RECT 0.146 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.37 0.194 ;
        RECT 0.274 0.638 0.37 0.666 ;
        RECT 0.37 0.166 0.398 0.194 ;
        RECT 0.37 0.194 0.398 0.376 ;
        RECT 0.37 0.376 0.398 0.638 ;
        RECT 0.37 0.638 0.398 0.666 ;
        RECT 0.398 0.638 0.56 0.666 ;
        RECT 0.56 0.376 0.588 0.638 ;
        RECT 0.56 0.638 0.588 0.666 ;
      LAYER M1 ;
        RECT 0.05 0.072 0.078 0.312 ;
        RECT 0.05 0.312 0.078 0.34 ;
        RECT 0.05 0.34 0.078 0.418 ;
        RECT 0.05 0.418 0.078 0.686 ;
        RECT 0.078 0.312 0.178 0.34 ;
        RECT 0.178 0.312 0.206 0.34 ;
        RECT 0.178 0.34 0.206 0.418 ;
        RECT 0.146 0.574 0.202 0.602 ;
        RECT 0.202 0.1019 0.23 0.13 ;
        RECT 0.202 0.13 0.23 0.23 ;
        RECT 0.202 0.23 0.23 0.258 ;
        RECT 0.202 0.574 0.23 0.602 ;
        RECT 0.23 0.1019 0.306 0.13 ;
        RECT 0.23 0.23 0.306 0.258 ;
        RECT 0.23 0.574 0.306 0.602 ;
        RECT 0.306 0.1019 0.334 0.13 ;
        RECT 0.306 0.23 0.334 0.258 ;
        RECT 0.306 0.258 0.334 0.314 ;
        RECT 0.306 0.314 0.334 0.574 ;
        RECT 0.306 0.574 0.334 0.602 ;
        RECT 0.334 0.1019 0.51 0.13 ;
        RECT 0.51 0.1019 0.542 0.13 ;
        RECT 0.51 0.13 0.542 0.23 ;
        RECT 0.51 0.23 0.542 0.258 ;
        RECT 0.51 0.258 0.542 0.314 ;
        RECT 0.146 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.37 0.194 ;
        RECT 0.274 0.638 0.37 0.666 ;
        RECT 0.37 0.166 0.398 0.194 ;
        RECT 0.37 0.194 0.398 0.376 ;
        RECT 0.37 0.376 0.398 0.638 ;
        RECT 0.37 0.638 0.398 0.666 ;
        RECT 0.398 0.638 0.56 0.666 ;
        RECT 0.56 0.376 0.588 0.638 ;
        RECT 0.56 0.638 0.588 0.666 ;
  END
END TBUF_X1

MACRO TBUF_X2
  CLASS core ;
  FOREIGN TBUF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.768 BY 0.768 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.384 0.1419 0.504 ;
        RECT 0.114 0.504 0.1419 0.532 ;
        RECT 0.1419 0.504 0.206 0.532 ;
        RECT 0.206 0.504 0.242 0.532 ;
        RECT 0.242 0.306 0.27 0.384 ;
        RECT 0.242 0.384 0.27 0.504 ;
        RECT 0.242 0.504 0.27 0.532 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.382 0.462 0.576 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.624 0.07 0.656 0.6959 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.53 0.796 ;
        RECT 0.53 0.74 0.778 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.778 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.072 0.078 0.312 ;
        RECT 0.05 0.312 0.078 0.34 ;
        RECT 0.05 0.34 0.078 0.404 ;
        RECT 0.05 0.404 0.078 0.612 ;
        RECT 0.078 0.312 0.178 0.34 ;
        RECT 0.178 0.312 0.206 0.34 ;
        RECT 0.178 0.34 0.206 0.404 ;
        RECT 0.146 0.5679 0.202 0.602 ;
        RECT 0.202 0.1019 0.23 0.13 ;
        RECT 0.202 0.13 0.23 0.23 ;
        RECT 0.202 0.23 0.23 0.258 ;
        RECT 0.202 0.5679 0.23 0.602 ;
        RECT 0.23 0.1019 0.306 0.13 ;
        RECT 0.23 0.23 0.306 0.258 ;
        RECT 0.23 0.5679 0.306 0.602 ;
        RECT 0.306 0.1019 0.334 0.13 ;
        RECT 0.306 0.23 0.334 0.258 ;
        RECT 0.306 0.258 0.334 0.314 ;
        RECT 0.306 0.314 0.334 0.5679 ;
        RECT 0.306 0.5679 0.334 0.602 ;
        RECT 0.334 0.1019 0.482 0.13 ;
        RECT 0.482 0.1019 0.514 0.13 ;
        RECT 0.482 0.13 0.514 0.23 ;
        RECT 0.482 0.23 0.514 0.258 ;
        RECT 0.482 0.258 0.514 0.314 ;
        RECT 0.146 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.37 0.194 ;
        RECT 0.274 0.638 0.37 0.666 ;
        RECT 0.37 0.166 0.398 0.194 ;
        RECT 0.37 0.194 0.398 0.443 ;
        RECT 0.37 0.443 0.398 0.638 ;
        RECT 0.37 0.638 0.398 0.666 ;
        RECT 0.398 0.638 0.498 0.666 ;
        RECT 0.498 0.443 0.53 0.638 ;
        RECT 0.498 0.638 0.53 0.666 ;
      LAYER M1 ;
        RECT 0.05 0.072 0.078 0.312 ;
        RECT 0.05 0.312 0.078 0.34 ;
        RECT 0.05 0.34 0.078 0.404 ;
        RECT 0.05 0.404 0.078 0.612 ;
        RECT 0.078 0.312 0.178 0.34 ;
        RECT 0.178 0.312 0.206 0.34 ;
        RECT 0.178 0.34 0.206 0.404 ;
        RECT 0.146 0.5679 0.202 0.602 ;
        RECT 0.202 0.1019 0.23 0.13 ;
        RECT 0.202 0.13 0.23 0.23 ;
        RECT 0.202 0.23 0.23 0.258 ;
        RECT 0.202 0.5679 0.23 0.602 ;
        RECT 0.23 0.1019 0.306 0.13 ;
        RECT 0.23 0.23 0.306 0.258 ;
        RECT 0.23 0.5679 0.306 0.602 ;
        RECT 0.306 0.1019 0.334 0.13 ;
        RECT 0.306 0.23 0.334 0.258 ;
        RECT 0.306 0.258 0.334 0.314 ;
        RECT 0.306 0.314 0.334 0.5679 ;
        RECT 0.306 0.5679 0.334 0.602 ;
        RECT 0.334 0.1019 0.482 0.13 ;
        RECT 0.482 0.1019 0.514 0.13 ;
        RECT 0.482 0.13 0.514 0.23 ;
        RECT 0.482 0.23 0.514 0.258 ;
        RECT 0.482 0.258 0.514 0.314 ;
        RECT 0.146 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.37 0.194 ;
        RECT 0.274 0.638 0.37 0.666 ;
        RECT 0.37 0.166 0.398 0.194 ;
        RECT 0.37 0.194 0.398 0.443 ;
        RECT 0.37 0.443 0.398 0.638 ;
        RECT 0.37 0.638 0.398 0.666 ;
        RECT 0.398 0.638 0.498 0.666 ;
        RECT 0.498 0.443 0.53 0.638 ;
        RECT 0.498 0.638 0.53 0.666 ;
  END
END TBUF_X2

MACRO TBUF_X4
  CLASS core ;
  FOREIGN TBUF_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.96 BY 0.768 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.384 0.1419 0.484 ;
        RECT 0.114 0.484 0.1419 0.512 ;
        RECT 0.1419 0.484 0.206 0.512 ;
        RECT 0.206 0.484 0.242 0.512 ;
        RECT 0.242 0.306 0.27 0.384 ;
        RECT 0.242 0.384 0.27 0.484 ;
        RECT 0.242 0.484 0.27 0.512 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.3459 0.462 0.594 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.6879 0.064 0.72 0.224 ;
        RECT 0.6879 0.224 0.72 0.256 ;
        RECT 0.6879 0.512 0.72 0.54 ;
        RECT 0.6879 0.54 0.72 0.5709 ;
        RECT 0.6879 0.5709 0.72 0.704 ;
        RECT 0.72 0.224 0.8129 0.256 ;
        RECT 0.72 0.512 0.8129 0.54 ;
        RECT 0.8129 0.064 0.8139 0.224 ;
        RECT 0.8129 0.224 0.8139 0.256 ;
        RECT 0.8129 0.512 0.8139 0.54 ;
        RECT 0.8139 0.064 0.8159 0.224 ;
        RECT 0.8139 0.224 0.8159 0.256 ;
        RECT 0.8139 0.512 0.8159 0.54 ;
        RECT 0.8159 0.064 0.838 0.224 ;
        RECT 0.8159 0.224 0.838 0.256 ;
        RECT 0.8159 0.512 0.838 0.54 ;
        RECT 0.8159 0.54 0.838 0.5709 ;
        RECT 0.8159 0.5709 0.838 0.704 ;
        RECT 0.838 0.064 0.848 0.224 ;
        RECT 0.838 0.224 0.848 0.256 ;
        RECT 0.838 0.512 0.848 0.54 ;
        RECT 0.838 0.54 0.848 0.5709 ;
        RECT 0.838 0.5709 0.848 0.704 ;
        RECT 0.848 0.064 0.851 0.224 ;
        RECT 0.848 0.224 0.851 0.256 ;
        RECT 0.848 0.512 0.851 0.54 ;
        RECT 0.848 0.54 0.851 0.5709 ;
        RECT 0.851 0.224 0.882 0.256 ;
        RECT 0.851 0.512 0.882 0.54 ;
        RECT 0.851 0.54 0.882 0.5709 ;
        RECT 0.882 0.224 0.91 0.256 ;
        RECT 0.882 0.256 0.91 0.512 ;
        RECT 0.882 0.512 0.91 0.54 ;
        RECT 0.882 0.54 0.91 0.5709 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.8139 0.796 ;
        RECT 0.8139 0.74 0.838 0.796 ;
        RECT 0.838 0.74 0.97 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.97 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.082 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.37 0.194 ;
        RECT 0.274 0.638 0.37 0.666 ;
        RECT 0.37 0.166 0.398 0.194 ;
        RECT 0.37 0.194 0.398 0.388 ;
        RECT 0.37 0.388 0.398 0.414 ;
        RECT 0.37 0.414 0.398 0.458 ;
        RECT 0.37 0.458 0.398 0.638 ;
        RECT 0.37 0.638 0.398 0.666 ;
        RECT 0.398 0.638 0.526 0.666 ;
        RECT 0.526 0.388 0.582 0.414 ;
        RECT 0.526 0.414 0.582 0.458 ;
        RECT 0.526 0.458 0.582 0.638 ;
        RECT 0.526 0.638 0.582 0.666 ;
        RECT 0.582 0.414 0.8139 0.458 ;
        RECT 0.05 0.096 0.078 0.312 ;
        RECT 0.05 0.312 0.078 0.34 ;
        RECT 0.05 0.34 0.078 0.404 ;
        RECT 0.05 0.404 0.078 0.594 ;
        RECT 0.078 0.312 0.178 0.34 ;
        RECT 0.178 0.312 0.206 0.34 ;
        RECT 0.178 0.34 0.206 0.404 ;
        RECT 0.146 0.5679 0.202 0.602 ;
        RECT 0.202 0.1019 0.23 0.13 ;
        RECT 0.202 0.13 0.23 0.23 ;
        RECT 0.202 0.23 0.23 0.258 ;
        RECT 0.202 0.5679 0.23 0.602 ;
        RECT 0.23 0.1019 0.306 0.13 ;
        RECT 0.23 0.23 0.306 0.258 ;
        RECT 0.23 0.5679 0.306 0.602 ;
        RECT 0.306 0.1019 0.334 0.13 ;
        RECT 0.306 0.23 0.334 0.258 ;
        RECT 0.306 0.258 0.334 0.292 ;
        RECT 0.306 0.292 0.334 0.32 ;
        RECT 0.306 0.32 0.334 0.352 ;
        RECT 0.306 0.352 0.334 0.5679 ;
        RECT 0.306 0.5679 0.334 0.602 ;
        RECT 0.334 0.1019 0.526 0.13 ;
        RECT 0.526 0.1019 0.582 0.13 ;
        RECT 0.526 0.13 0.582 0.23 ;
        RECT 0.526 0.23 0.582 0.258 ;
        RECT 0.526 0.258 0.582 0.292 ;
        RECT 0.526 0.292 0.582 0.32 ;
        RECT 0.526 0.32 0.582 0.352 ;
        RECT 0.582 0.292 0.838 0.32 ;
      LAYER M1 ;
        RECT 0.082 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.37 0.194 ;
        RECT 0.274 0.638 0.37 0.666 ;
        RECT 0.37 0.166 0.398 0.194 ;
        RECT 0.37 0.194 0.398 0.388 ;
        RECT 0.37 0.388 0.398 0.414 ;
        RECT 0.37 0.414 0.398 0.458 ;
        RECT 0.37 0.458 0.398 0.638 ;
        RECT 0.37 0.638 0.398 0.666 ;
        RECT 0.398 0.638 0.526 0.666 ;
        RECT 0.526 0.388 0.582 0.414 ;
        RECT 0.526 0.414 0.582 0.458 ;
        RECT 0.526 0.458 0.582 0.638 ;
        RECT 0.526 0.638 0.582 0.666 ;
        RECT 0.582 0.414 0.8139 0.458 ;
        RECT 0.05 0.096 0.078 0.312 ;
        RECT 0.05 0.312 0.078 0.34 ;
        RECT 0.05 0.34 0.078 0.404 ;
        RECT 0.05 0.404 0.078 0.594 ;
        RECT 0.078 0.312 0.178 0.34 ;
        RECT 0.178 0.312 0.206 0.34 ;
        RECT 0.178 0.34 0.206 0.404 ;
        RECT 0.146 0.5679 0.202 0.602 ;
        RECT 0.202 0.1019 0.23 0.13 ;
        RECT 0.202 0.13 0.23 0.23 ;
        RECT 0.202 0.23 0.23 0.258 ;
        RECT 0.202 0.5679 0.23 0.602 ;
        RECT 0.23 0.1019 0.306 0.13 ;
        RECT 0.23 0.23 0.306 0.258 ;
        RECT 0.23 0.5679 0.306 0.602 ;
        RECT 0.306 0.1019 0.334 0.13 ;
        RECT 0.306 0.23 0.334 0.258 ;
        RECT 0.306 0.258 0.334 0.292 ;
        RECT 0.306 0.292 0.334 0.32 ;
        RECT 0.306 0.32 0.334 0.352 ;
        RECT 0.306 0.352 0.334 0.5679 ;
        RECT 0.306 0.5679 0.334 0.602 ;
        RECT 0.334 0.1019 0.526 0.13 ;
        RECT 0.526 0.1019 0.582 0.13 ;
        RECT 0.526 0.13 0.582 0.23 ;
        RECT 0.526 0.23 0.582 0.258 ;
        RECT 0.526 0.258 0.582 0.292 ;
        RECT 0.526 0.292 0.582 0.32 ;
        RECT 0.526 0.32 0.582 0.352 ;
        RECT 0.582 0.292 0.838 0.32 ;
  END
END TBUF_X4

MACRO TBUF_X8
  CLASS core ;
  FOREIGN TBUF_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.344 BY 0.768 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.384 0.1419 0.484 ;
        RECT 0.114 0.484 0.1419 0.512 ;
        RECT 0.1419 0.484 0.222 0.512 ;
        RECT 0.222 0.484 0.306 0.512 ;
        RECT 0.306 0.32 0.334 0.384 ;
        RECT 0.306 0.384 0.334 0.484 ;
        RECT 0.306 0.484 0.334 0.512 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.498 0.3459 0.526 0.402 ;
        RECT 0.498 0.402 0.526 0.434 ;
        RECT 0.498 0.434 0.526 0.576 ;
        RECT 0.526 0.402 0.622 0.434 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.8159 0.064 0.848 0.133 ;
        RECT 0.8159 0.133 0.848 0.16 ;
        RECT 0.8159 0.16 0.848 0.192 ;
        RECT 0.8159 0.519 0.848 0.577 ;
        RECT 0.8159 0.577 0.848 0.578 ;
        RECT 0.8159 0.578 0.848 0.704 ;
        RECT 0.848 0.16 1.183 0.192 ;
        RECT 0.848 0.519 1.183 0.577 ;
        RECT 1.183 0.16 1.198 0.192 ;
        RECT 1.183 0.519 1.198 0.577 ;
        RECT 1.198 0.16 1.2 0.192 ;
        RECT 1.198 0.519 1.2 0.577 ;
        RECT 1.2 0.064 1.232 0.133 ;
        RECT 1.2 0.133 1.232 0.16 ;
        RECT 1.2 0.16 1.232 0.192 ;
        RECT 1.2 0.519 1.232 0.577 ;
        RECT 1.2 0.577 1.232 0.578 ;
        RECT 1.2 0.578 1.232 0.704 ;
        RECT 1.232 0.133 1.266 0.16 ;
        RECT 1.232 0.16 1.266 0.192 ;
        RECT 1.232 0.519 1.266 0.577 ;
        RECT 1.232 0.577 1.266 0.578 ;
        RECT 1.266 0.133 1.294 0.16 ;
        RECT 1.266 0.16 1.294 0.192 ;
        RECT 1.266 0.192 1.294 0.519 ;
        RECT 1.266 0.519 1.294 0.577 ;
        RECT 1.266 0.577 1.294 0.578 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.183 0.796 ;
        RECT 1.183 0.74 1.198 0.796 ;
        RECT 1.198 0.74 1.354 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.354 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.072 0.078 0.312 ;
        RECT 0.05 0.312 0.078 0.34 ;
        RECT 0.05 0.34 0.078 0.43 ;
        RECT 0.05 0.43 0.078 0.638 ;
        RECT 0.078 0.312 0.178 0.34 ;
        RECT 0.178 0.312 0.222 0.34 ;
        RECT 0.178 0.34 0.222 0.43 ;
        RECT 0.146 0.574 0.202 0.602 ;
        RECT 0.202 0.1019 0.23 0.13 ;
        RECT 0.202 0.13 0.23 0.23 ;
        RECT 0.202 0.23 0.23 0.258 ;
        RECT 0.202 0.574 0.23 0.602 ;
        RECT 0.23 0.1019 0.37 0.13 ;
        RECT 0.23 0.23 0.37 0.258 ;
        RECT 0.23 0.574 0.37 0.602 ;
        RECT 0.37 0.1019 0.398 0.13 ;
        RECT 0.37 0.23 0.398 0.258 ;
        RECT 0.37 0.258 0.398 0.2859 ;
        RECT 0.37 0.2859 0.398 0.342 ;
        RECT 0.37 0.342 0.398 0.574 ;
        RECT 0.37 0.574 0.398 0.602 ;
        RECT 0.398 0.1019 0.6899 0.13 ;
        RECT 0.6899 0.1019 0.718 0.13 ;
        RECT 0.6899 0.13 0.718 0.23 ;
        RECT 0.6899 0.23 0.718 0.258 ;
        RECT 0.6899 0.258 0.718 0.2859 ;
        RECT 0.6899 0.2859 0.718 0.342 ;
        RECT 0.718 0.258 1.198 0.2859 ;
        RECT 0.122 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.434 0.194 ;
        RECT 0.274 0.638 0.434 0.666 ;
        RECT 0.434 0.166 0.462 0.194 ;
        RECT 0.434 0.194 0.462 0.386 ;
        RECT 0.434 0.386 0.462 0.403 ;
        RECT 0.434 0.403 0.462 0.461 ;
        RECT 0.434 0.461 0.462 0.638 ;
        RECT 0.434 0.638 0.462 0.666 ;
        RECT 0.462 0.638 0.66 0.666 ;
        RECT 0.66 0.386 0.718 0.403 ;
        RECT 0.66 0.403 0.718 0.461 ;
        RECT 0.66 0.461 0.718 0.638 ;
        RECT 0.66 0.638 0.718 0.666 ;
        RECT 0.718 0.403 1.183 0.461 ;
      LAYER M1 ;
        RECT 0.05 0.072 0.078 0.312 ;
        RECT 0.05 0.312 0.078 0.34 ;
        RECT 0.05 0.34 0.078 0.43 ;
        RECT 0.05 0.43 0.078 0.638 ;
        RECT 0.078 0.312 0.178 0.34 ;
        RECT 0.178 0.312 0.222 0.34 ;
        RECT 0.178 0.34 0.222 0.43 ;
        RECT 0.146 0.574 0.202 0.602 ;
        RECT 0.202 0.1019 0.23 0.13 ;
        RECT 0.202 0.13 0.23 0.23 ;
        RECT 0.202 0.23 0.23 0.258 ;
        RECT 0.202 0.574 0.23 0.602 ;
        RECT 0.23 0.1019 0.37 0.13 ;
        RECT 0.23 0.23 0.37 0.258 ;
        RECT 0.23 0.574 0.37 0.602 ;
        RECT 0.37 0.1019 0.398 0.13 ;
        RECT 0.37 0.23 0.398 0.258 ;
        RECT 0.37 0.258 0.398 0.2859 ;
        RECT 0.37 0.2859 0.398 0.342 ;
        RECT 0.37 0.342 0.398 0.574 ;
        RECT 0.37 0.574 0.398 0.602 ;
        RECT 0.398 0.1019 0.6899 0.13 ;
        RECT 0.6899 0.1019 0.718 0.13 ;
        RECT 0.6899 0.13 0.718 0.23 ;
        RECT 0.6899 0.23 0.718 0.258 ;
        RECT 0.6899 0.258 0.718 0.2859 ;
        RECT 0.6899 0.2859 0.718 0.342 ;
        RECT 0.718 0.258 1.198 0.2859 ;
        RECT 0.122 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.434 0.194 ;
        RECT 0.274 0.638 0.434 0.666 ;
        RECT 0.434 0.166 0.462 0.194 ;
        RECT 0.434 0.194 0.462 0.386 ;
        RECT 0.434 0.386 0.462 0.403 ;
        RECT 0.434 0.403 0.462 0.461 ;
        RECT 0.434 0.461 0.462 0.638 ;
        RECT 0.434 0.638 0.462 0.666 ;
        RECT 0.462 0.638 0.66 0.666 ;
        RECT 0.66 0.386 0.718 0.403 ;
        RECT 0.66 0.403 0.718 0.461 ;
        RECT 0.66 0.461 0.718 0.638 ;
        RECT 0.66 0.638 0.718 0.666 ;
        RECT 0.718 0.403 1.183 0.461 ;
  END
END TBUF_X8

MACRO TBUF_X12
  CLASS core ;
  FOREIGN TBUF_X12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 1.728 BY 0.768 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.384 0.1419 0.51 ;
        RECT 0.114 0.51 0.1419 0.538 ;
        RECT 0.1419 0.51 0.206 0.538 ;
        RECT 0.206 0.51 0.242 0.538 ;
        RECT 0.242 0.306 0.27 0.384 ;
        RECT 0.242 0.384 0.27 0.51 ;
        RECT 0.242 0.51 0.27 0.538 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.434 0.402 0.498 0.448 ;
        RECT 0.498 0.3459 0.526 0.402 ;
        RECT 0.498 0.402 0.526 0.448 ;
        RECT 0.526 0.402 0.626 0.448 ;
        RECT 0.626 0.402 0.654 0.448 ;
        RECT 0.626 0.448 0.654 0.576 ;
        RECT 0.654 0.402 0.71 0.448 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.684 0.796 ;
        RECT 1.684 0.74 1.738 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 1.738 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.146 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.37 0.194 ;
        RECT 0.274 0.638 0.37 0.666 ;
        RECT 0.37 0.166 0.398 0.194 ;
        RECT 0.37 0.194 0.398 0.356 ;
        RECT 0.37 0.356 0.398 0.378 ;
        RECT 0.37 0.378 0.398 0.426 ;
        RECT 0.37 0.426 0.398 0.638 ;
        RECT 0.37 0.638 0.398 0.666 ;
        RECT 0.398 0.638 0.783 0.666 ;
        RECT 0.783 0.356 0.839 0.378 ;
        RECT 0.783 0.378 0.839 0.426 ;
        RECT 0.783 0.426 0.839 0.638 ;
        RECT 0.783 0.638 0.839 0.666 ;
        RECT 0.839 0.378 1.557 0.426 ;
        RECT 0.882 0.1019 0.931 0.13 ;
        RECT 0.931 0.1019 0.989 0.13 ;
        RECT 0.931 0.532 0.989 0.5639 ;
        RECT 0.931 0.5639 0.989 0.62 ;
        RECT 0.989 0.1019 1.572 0.13 ;
        RECT 0.989 0.532 1.572 0.5639 ;
        RECT 1.572 0.073 1.586 0.1019 ;
        RECT 1.572 0.1019 1.586 0.13 ;
        RECT 1.572 0.532 1.586 0.5639 ;
        RECT 1.586 0.073 1.614 0.1019 ;
        RECT 1.586 0.1019 1.614 0.13 ;
        RECT 1.586 0.532 1.614 0.5639 ;
        RECT 1.586 0.5639 1.614 0.62 ;
        RECT 1.586 0.62 1.614 0.624 ;
        RECT 1.614 0.073 1.6279 0.1019 ;
        RECT 1.614 0.1019 1.6279 0.13 ;
        RECT 1.614 0.532 1.6279 0.5639 ;
        RECT 1.6279 0.1019 1.629 0.13 ;
        RECT 1.6279 0.532 1.629 0.5639 ;
        RECT 1.629 0.1019 1.684 0.13 ;
        RECT 1.629 0.13 1.684 0.532 ;
        RECT 1.629 0.532 1.684 0.5639 ;
        RECT 0.05 0.1739 0.078 0.312 ;
        RECT 0.05 0.312 0.078 0.34 ;
        RECT 0.05 0.34 0.078 0.404 ;
        RECT 0.05 0.404 0.078 0.672 ;
        RECT 0.078 0.312 0.178 0.34 ;
        RECT 0.178 0.312 0.206 0.34 ;
        RECT 0.178 0.34 0.206 0.404 ;
        RECT 0.1419 0.1019 0.146 0.13 ;
        RECT 0.1419 0.13 0.146 0.23 ;
        RECT 0.1419 0.23 0.146 0.25 ;
        RECT 0.1419 0.25 0.146 0.258 ;
        RECT 0.146 0.1019 0.17 0.13 ;
        RECT 0.146 0.13 0.17 0.23 ;
        RECT 0.146 0.23 0.17 0.25 ;
        RECT 0.146 0.25 0.17 0.258 ;
        RECT 0.146 0.574 0.17 0.602 ;
        RECT 0.17 0.1019 0.306 0.13 ;
        RECT 0.17 0.23 0.306 0.25 ;
        RECT 0.17 0.25 0.306 0.258 ;
        RECT 0.17 0.574 0.306 0.602 ;
        RECT 0.306 0.1019 0.334 0.13 ;
        RECT 0.306 0.23 0.334 0.25 ;
        RECT 0.306 0.25 0.334 0.258 ;
        RECT 0.306 0.258 0.334 0.294 ;
        RECT 0.306 0.294 0.334 0.574 ;
        RECT 0.306 0.574 0.334 0.602 ;
        RECT 0.334 0.1019 0.782 0.13 ;
        RECT 0.782 0.1019 0.8139 0.13 ;
        RECT 0.782 0.13 0.8139 0.23 ;
        RECT 0.782 0.23 0.8139 0.25 ;
        RECT 0.782 0.25 0.8139 0.258 ;
        RECT 0.782 0.258 0.8139 0.294 ;
        RECT 0.8139 0.25 1.593 0.258 ;
        RECT 0.8139 0.258 1.593 0.294 ;
      LAYER M1 ;
        RECT 0.146 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.37 0.194 ;
        RECT 0.274 0.638 0.37 0.666 ;
        RECT 0.37 0.166 0.398 0.194 ;
        RECT 0.37 0.194 0.398 0.356 ;
        RECT 0.37 0.356 0.398 0.378 ;
        RECT 0.37 0.378 0.398 0.426 ;
        RECT 0.37 0.426 0.398 0.638 ;
        RECT 0.37 0.638 0.398 0.666 ;
        RECT 0.398 0.638 0.783 0.666 ;
        RECT 0.783 0.356 0.839 0.378 ;
        RECT 0.783 0.378 0.839 0.426 ;
        RECT 0.783 0.426 0.839 0.638 ;
        RECT 0.783 0.638 0.839 0.666 ;
        RECT 0.839 0.378 1.557 0.426 ;
        RECT 0.882 0.1019 0.931 0.13 ;
        RECT 0.931 0.1019 0.989 0.13 ;
        RECT 0.931 0.532 0.989 0.5639 ;
        RECT 0.931 0.5639 0.989 0.62 ;
        RECT 0.989 0.1019 1.572 0.13 ;
        RECT 0.989 0.532 1.572 0.5639 ;
        RECT 1.572 0.073 1.586 0.1019 ;
        RECT 1.572 0.1019 1.586 0.13 ;
        RECT 1.572 0.532 1.586 0.5639 ;
        RECT 1.586 0.073 1.614 0.1019 ;
        RECT 1.586 0.1019 1.614 0.13 ;
        RECT 1.586 0.532 1.614 0.5639 ;
        RECT 1.586 0.5639 1.614 0.62 ;
        RECT 1.586 0.62 1.614 0.624 ;
        RECT 1.614 0.073 1.6279 0.1019 ;
        RECT 1.614 0.1019 1.6279 0.13 ;
        RECT 1.614 0.532 1.6279 0.5639 ;
        RECT 1.6279 0.1019 1.629 0.13 ;
        RECT 1.6279 0.532 1.629 0.5639 ;
        RECT 1.629 0.1019 1.684 0.13 ;
        RECT 1.629 0.13 1.684 0.532 ;
        RECT 1.629 0.532 1.684 0.5639 ;
        RECT 0.05 0.1739 0.078 0.312 ;
        RECT 0.05 0.312 0.078 0.34 ;
        RECT 0.05 0.34 0.078 0.404 ;
        RECT 0.05 0.404 0.078 0.672 ;
        RECT 0.078 0.312 0.178 0.34 ;
        RECT 0.178 0.312 0.206 0.34 ;
        RECT 0.178 0.34 0.206 0.404 ;
        RECT 0.1419 0.1019 0.146 0.13 ;
        RECT 0.1419 0.13 0.146 0.23 ;
        RECT 0.1419 0.23 0.146 0.25 ;
        RECT 0.1419 0.25 0.146 0.258 ;
        RECT 0.146 0.1019 0.17 0.13 ;
        RECT 0.146 0.13 0.17 0.23 ;
        RECT 0.146 0.23 0.17 0.25 ;
        RECT 0.146 0.25 0.17 0.258 ;
        RECT 0.146 0.574 0.17 0.602 ;
        RECT 0.17 0.1019 0.306 0.13 ;
        RECT 0.17 0.23 0.306 0.25 ;
        RECT 0.17 0.25 0.306 0.258 ;
        RECT 0.17 0.574 0.306 0.602 ;
        RECT 0.306 0.1019 0.334 0.13 ;
        RECT 0.306 0.23 0.334 0.25 ;
        RECT 0.306 0.25 0.334 0.258 ;
        RECT 0.306 0.258 0.334 0.294 ;
        RECT 0.306 0.294 0.334 0.574 ;
        RECT 0.306 0.574 0.334 0.602 ;
        RECT 0.334 0.1019 0.782 0.13 ;
        RECT 0.782 0.1019 0.8139 0.13 ;
        RECT 0.782 0.13 0.8139 0.23 ;
        RECT 0.782 0.23 0.8139 0.25 ;
        RECT 0.782 0.25 0.8139 0.258 ;
        RECT 0.782 0.258 0.8139 0.294 ;
        RECT 0.8139 0.25 1.593 0.258 ;
        RECT 0.8139 0.258 1.593 0.294 ;
  END
END TBUF_X12

MACRO TBUF_X16
  CLASS core ;
  FOREIGN TBUF_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 2.112 BY 0.768 ;
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.114 0.39 0.1419 0.486 ;
        RECT 0.114 0.486 0.1419 0.514 ;
        RECT 0.1419 0.486 0.1739 0.514 ;
        RECT 0.1739 0.486 0.24 0.514 ;
        RECT 0.24 0.32 0.272 0.39 ;
        RECT 0.24 0.39 0.272 0.486 ;
        RECT 0.24 0.486 0.272 0.514 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.462 0.402 0.562 0.448 ;
        RECT 0.562 0.3459 0.59 0.402 ;
        RECT 0.562 0.402 0.59 0.448 ;
        RECT 0.59 0.402 0.6899 0.448 ;
        RECT 0.6899 0.402 0.718 0.448 ;
        RECT 0.6899 0.448 0.718 0.576 ;
        RECT 0.718 0.402 0.902 0.448 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 1.072 0.064 1.104 0.1419 ;
        RECT 1.072 0.1419 1.104 0.2 ;
        RECT 1.072 0.52 1.104 0.576 ;
        RECT 1.072 0.576 1.104 0.704 ;
        RECT 1.104 0.1419 1.968 0.2 ;
        RECT 1.104 0.52 1.968 0.576 ;
        RECT 1.968 0.064 1.98 0.1419 ;
        RECT 1.968 0.1419 1.98 0.2 ;
        RECT 1.968 0.52 1.98 0.576 ;
        RECT 1.968 0.576 1.98 0.704 ;
        RECT 1.98 0.064 1.998 0.1419 ;
        RECT 1.98 0.1419 1.998 0.2 ;
        RECT 1.98 0.52 1.998 0.576 ;
        RECT 1.98 0.576 1.998 0.704 ;
        RECT 1.998 0.064 2 0.1419 ;
        RECT 1.998 0.1419 2 0.2 ;
        RECT 1.998 0.52 2 0.576 ;
        RECT 1.998 0.576 2 0.704 ;
        RECT 2 0.1419 2.0339 0.2 ;
        RECT 2 0.52 2.0339 0.576 ;
        RECT 2.0339 0.1419 2.062 0.2 ;
        RECT 2.0339 0.2 2.062 0.52 ;
        RECT 2.0339 0.52 2.062 0.576 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 1.98 0.796 ;
        RECT 1.98 0.74 1.998 0.796 ;
        RECT 1.998 0.74 2.122 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 2.122 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.05 0.072 0.078 0.262 ;
        RECT 0.05 0.262 0.078 0.29 ;
        RECT 0.05 0.29 0.078 0.3459 ;
        RECT 0.05 0.3459 0.078 0.6 ;
        RECT 0.078 0.262 0.1419 0.29 ;
        RECT 0.1419 0.262 0.1739 0.29 ;
        RECT 0.1419 0.29 0.1739 0.3459 ;
        RECT 0.146 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.398 0.198 ;
        RECT 0.274 0.638 0.398 0.666 ;
        RECT 0.398 0.166 0.426 0.198 ;
        RECT 0.398 0.198 0.426 0.403 ;
        RECT 0.398 0.403 0.426 0.461 ;
        RECT 0.398 0.461 0.426 0.638 ;
        RECT 0.398 0.638 0.426 0.666 ;
        RECT 0.426 0.638 0.946 0.666 ;
        RECT 0.946 0.403 0.974 0.461 ;
        RECT 0.946 0.461 0.974 0.638 ;
        RECT 0.946 0.638 0.974 0.666 ;
        RECT 0.974 0.403 1.98 0.461 ;
        RECT 0.146 0.5679 0.21 0.602 ;
        RECT 0.21 0.1019 0.238 0.13 ;
        RECT 0.21 0.13 0.238 0.234 ;
        RECT 0.21 0.234 0.238 0.262 ;
        RECT 0.21 0.5679 0.238 0.602 ;
        RECT 0.238 0.1019 0.326 0.13 ;
        RECT 0.238 0.234 0.326 0.262 ;
        RECT 0.238 0.5679 0.326 0.602 ;
        RECT 0.326 0.1019 0.362 0.13 ;
        RECT 0.326 0.234 0.362 0.262 ;
        RECT 0.326 0.262 0.362 0.273 ;
        RECT 0.326 0.273 0.362 0.331 ;
        RECT 0.326 0.331 0.362 0.5679 ;
        RECT 0.326 0.5679 0.362 0.602 ;
        RECT 0.362 0.1019 0.946 0.13 ;
        RECT 0.946 0.1019 0.974 0.13 ;
        RECT 0.946 0.13 0.974 0.234 ;
        RECT 0.946 0.234 0.974 0.262 ;
        RECT 0.946 0.262 0.974 0.273 ;
        RECT 0.946 0.273 0.974 0.331 ;
        RECT 0.974 0.273 1.998 0.331 ;
      LAYER M1 ;
        RECT 0.05 0.072 0.078 0.262 ;
        RECT 0.05 0.262 0.078 0.29 ;
        RECT 0.05 0.29 0.078 0.3459 ;
        RECT 0.05 0.3459 0.078 0.6 ;
        RECT 0.078 0.262 0.1419 0.29 ;
        RECT 0.1419 0.262 0.1739 0.29 ;
        RECT 0.1419 0.29 0.1739 0.3459 ;
        RECT 0.146 0.638 0.274 0.666 ;
        RECT 0.274 0.166 0.398 0.198 ;
        RECT 0.274 0.638 0.398 0.666 ;
        RECT 0.398 0.166 0.426 0.198 ;
        RECT 0.398 0.198 0.426 0.403 ;
        RECT 0.398 0.403 0.426 0.461 ;
        RECT 0.398 0.461 0.426 0.638 ;
        RECT 0.398 0.638 0.426 0.666 ;
        RECT 0.426 0.638 0.946 0.666 ;
        RECT 0.946 0.403 0.974 0.461 ;
        RECT 0.946 0.461 0.974 0.638 ;
        RECT 0.946 0.638 0.974 0.666 ;
        RECT 0.974 0.403 1.98 0.461 ;
        RECT 0.146 0.5679 0.21 0.602 ;
        RECT 0.21 0.1019 0.238 0.13 ;
        RECT 0.21 0.13 0.238 0.234 ;
        RECT 0.21 0.234 0.238 0.262 ;
        RECT 0.21 0.5679 0.238 0.602 ;
        RECT 0.238 0.1019 0.326 0.13 ;
        RECT 0.238 0.234 0.326 0.262 ;
        RECT 0.238 0.5679 0.326 0.602 ;
        RECT 0.326 0.1019 0.362 0.13 ;
        RECT 0.326 0.234 0.362 0.262 ;
        RECT 0.326 0.262 0.362 0.273 ;
        RECT 0.326 0.273 0.362 0.331 ;
        RECT 0.326 0.331 0.362 0.5679 ;
        RECT 0.326 0.5679 0.362 0.602 ;
        RECT 0.362 0.1019 0.946 0.13 ;
        RECT 0.946 0.1019 0.974 0.13 ;
        RECT 0.946 0.13 0.974 0.234 ;
        RECT 0.946 0.234 0.974 0.262 ;
        RECT 0.946 0.262 0.974 0.273 ;
        RECT 0.946 0.273 0.974 0.331 ;
        RECT 0.974 0.273 1.998 0.331 ;
  END
END TBUF_X16

MACRO TIEH
  CLASS core ;
  FOREIGN TIEH 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.192 BY 0.768 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.109 0.473 0.1419 0.704 ;
        RECT 0.1419 0.473 0.147 0.704 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.1419 0.796 ;
        RECT 0.1419 0.74 0.202 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.202 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.096 0.1419 0.429 ;
      LAYER M1 ;
        RECT 0.114 0.096 0.1419 0.429 ;
  END
END TIEH

MACRO TIEL
  CLASS core ;
  FOREIGN TIEL 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.192 BY 0.768 ;
  PIN Z
    DIRECTION INOUT ;
    PORT
      LAYER M1 ;
        RECT 0.109 0.064 0.147 0.266 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.1419 0.796 ;
        RECT 0.1419 0.74 0.202 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.202 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.114 0.336 0.1419 0.672 ;
      LAYER M1 ;
        RECT 0.114 0.336 0.1419 0.672 ;
  END
END TIEL

MACRO XNOR2_X1
  CLASS core ;
  FOREIGN XNOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.252 0.21 0.28 ;
        RECT 0.178 0.28 0.21 0.428 ;
        RECT 0.21 0.252 0.37 0.28 ;
        RECT 0.37 0.252 0.398 0.28 ;
        RECT 0.37 0.28 0.398 0.428 ;
        RECT 0.37 0.428 0.398 0.448 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.242 0.078 0.32 ;
        RECT 0.05 0.32 0.078 0.676 ;
        RECT 0.05 0.676 0.078 0.704 ;
        RECT 0.078 0.676 0.274 0.704 ;
        RECT 0.274 0.676 0.498 0.704 ;
        RECT 0.498 0.32 0.526 0.676 ;
        RECT 0.498 0.676 0.526 0.704 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.278 0.546 0.302 0.547 ;
        RECT 0.278 0.547 0.302 0.601 ;
        RECT 0.278 0.601 0.302 0.602 ;
        RECT 0.302 0.166 0.334 0.194 ;
        RECT 0.302 0.546 0.334 0.547 ;
        RECT 0.302 0.547 0.334 0.601 ;
        RECT 0.302 0.601 0.334 0.602 ;
        RECT 0.334 0.166 0.434 0.194 ;
        RECT 0.334 0.547 0.434 0.601 ;
        RECT 0.434 0.166 0.462 0.194 ;
        RECT 0.434 0.248 0.462 0.276 ;
        RECT 0.434 0.276 0.462 0.546 ;
        RECT 0.434 0.546 0.462 0.547 ;
        RECT 0.434 0.547 0.462 0.601 ;
        RECT 0.462 0.166 0.493 0.194 ;
        RECT 0.462 0.248 0.493 0.276 ;
        RECT 0.493 0.166 0.531 0.194 ;
        RECT 0.493 0.194 0.531 0.248 ;
        RECT 0.493 0.248 0.531 0.276 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.274 0.796 ;
        RECT 0.274 0.74 0.535 0.796 ;
        RECT 0.535 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.21 0.1019 0.535 0.13 ;
        RECT 0.114 0.184 0.1419 0.216 ;
        RECT 0.114 0.216 0.1419 0.34 ;
        RECT 0.114 0.34 0.1419 0.464 ;
        RECT 0.114 0.464 0.1419 0.492 ;
        RECT 0.114 0.492 0.1419 0.552 ;
        RECT 0.1419 0.184 0.234 0.216 ;
        RECT 0.1419 0.464 0.234 0.492 ;
        RECT 0.234 0.464 0.246 0.492 ;
        RECT 0.246 0.34 0.274 0.464 ;
        RECT 0.246 0.464 0.274 0.492 ;
      LAYER M1 ;
        RECT 0.21 0.1019 0.535 0.13 ;
        RECT 0.114 0.184 0.1419 0.216 ;
        RECT 0.114 0.216 0.1419 0.34 ;
        RECT 0.114 0.34 0.1419 0.464 ;
        RECT 0.114 0.464 0.1419 0.492 ;
        RECT 0.114 0.492 0.1419 0.552 ;
        RECT 0.1419 0.184 0.234 0.216 ;
        RECT 0.1419 0.464 0.234 0.492 ;
        RECT 0.234 0.464 0.246 0.492 ;
        RECT 0.246 0.34 0.274 0.464 ;
        RECT 0.246 0.464 0.274 0.492 ;
  END
END XNOR2_X1

MACRO XOR2_X1
  CLASS core ;
  FOREIGN XOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NanGate_15nm_OCL ;
  SIZE 0.576 BY 0.768 ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.178 0.3439 0.21 0.486 ;
        RECT 0.178 0.486 0.21 0.514 ;
        RECT 0.21 0.486 0.274 0.514 ;
        RECT 0.274 0.486 0.37 0.514 ;
        RECT 0.37 0.32 0.398 0.3439 ;
        RECT 0.37 0.3439 0.398 0.486 ;
        RECT 0.37 0.486 0.398 0.514 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        RECT 0.05 0.064 0.078 0.092 ;
        RECT 0.05 0.092 0.078 0.448 ;
        RECT 0.05 0.448 0.078 0.526 ;
        RECT 0.078 0.064 0.498 0.092 ;
        RECT 0.498 0.064 0.526 0.092 ;
        RECT 0.498 0.092 0.526 0.448 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        RECT 0.275 0.163 0.315 0.164 ;
        RECT 0.275 0.164 0.315 0.222 ;
        RECT 0.315 0.163 0.334 0.164 ;
        RECT 0.315 0.164 0.334 0.222 ;
        RECT 0.315 0.574 0.334 0.602 ;
        RECT 0.334 0.164 0.434 0.222 ;
        RECT 0.334 0.574 0.434 0.602 ;
        RECT 0.434 0.164 0.462 0.222 ;
        RECT 0.434 0.222 0.462 0.492 ;
        RECT 0.434 0.492 0.462 0.52 ;
        RECT 0.434 0.574 0.462 0.602 ;
        RECT 0.462 0.492 0.496 0.52 ;
        RECT 0.462 0.574 0.496 0.602 ;
        RECT 0.496 0.492 0.528 0.52 ;
        RECT 0.496 0.52 0.528 0.574 ;
        RECT 0.496 0.574 0.528 0.602 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 0.74 0.535 0.796 ;
        RECT 0.535 0.74 0.586 0.796 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT -0.01 -0.028 0.586 0.028 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.246 0.638 0.535 0.666 ;
        RECT 0.114 0.136 0.1419 0.28 ;
        RECT 0.114 0.28 0.1419 0.308 ;
        RECT 0.114 0.308 0.1419 0.432 ;
        RECT 0.114 0.432 0.1419 0.552 ;
        RECT 0.114 0.552 0.1419 0.584 ;
        RECT 0.1419 0.28 0.246 0.308 ;
        RECT 0.1419 0.552 0.246 0.584 ;
        RECT 0.246 0.28 0.247 0.308 ;
        RECT 0.246 0.308 0.247 0.432 ;
        RECT 0.246 0.552 0.247 0.584 ;
        RECT 0.247 0.28 0.274 0.308 ;
        RECT 0.247 0.308 0.274 0.432 ;
      LAYER M1 ;
        RECT 0.246 0.638 0.535 0.666 ;
        RECT 0.114 0.136 0.1419 0.28 ;
        RECT 0.114 0.28 0.1419 0.308 ;
        RECT 0.114 0.308 0.1419 0.432 ;
        RECT 0.114 0.432 0.1419 0.552 ;
        RECT 0.114 0.552 0.1419 0.584 ;
        RECT 0.1419 0.28 0.246 0.308 ;
        RECT 0.1419 0.552 0.246 0.584 ;
        RECT 0.246 0.28 0.247 0.308 ;
        RECT 0.246 0.308 0.247 0.432 ;
        RECT 0.246 0.552 0.247 0.584 ;
        RECT 0.247 0.28 0.274 0.308 ;
        RECT 0.247 0.308 0.274 0.432 ;
  END
END XOR2_X1

END LIBRARY
#
# End of file
#
